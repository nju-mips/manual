`define RANDOMIZE_MEM_INIT
`define RANDOMIZE_REG_INIT
`define RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE_GARBAGE_ASSIGN
module RegFile(
  input         clock,
  input         reset,
  input         io_bp_valid,
  input         io_bp_bits_v,
  input  [4:0]  io_bp_bits_rd_idx,
  input         io_bp_bits_wen,
  input  [31:0] io_bp_bits_data,
  input         io_wb_valid,
  input         io_wb_bits_v,
  input  [7:0]  io_wb_bits_id,
  input  [31:0] io_wb_bits_pc,
  input  [5:0]  io_wb_bits_instr_op,
  input  [4:0]  io_wb_bits_instr_rs_idx,
  input  [4:0]  io_wb_bits_instr_rt_idx,
  input  [4:0]  io_wb_bits_instr_rd_idx,
  input  [4:0]  io_wb_bits_instr_shamt,
  input  [5:0]  io_wb_bits_instr_func,
  input  [4:0]  io_wb_bits_rd_idx,
  input         io_wb_bits_wen,
  input  [31:0] io_wb_bits_data,
  input         io_wb_bits_ip7,
  input  [4:0]  io_rfio_rs_idx,
  input  [4:0]  io_rfio_rt_idx,
  input         io_rfio_wen,
  input  [7:0]  io_rfio_wid,
  input  [4:0]  io_rfio_rd_idx,
  output        io_rfio_rs_data_valid,
  output [31:0] io_rfio_rs_data_bits,
  output        io_rfio_rt_data_valid,
  output [31:0] io_rfio_rt_data_bits,
  output        io_commit_valid,
  output [31:0] io_commit_pc,
  output [31:0] io_commit_instr,
  output        io_commit_ip7,
  output [31:0] io_commit_gpr_0,
  output [31:0] io_commit_gpr_1,
  output [31:0] io_commit_gpr_2,
  output [31:0] io_commit_gpr_3,
  output [31:0] io_commit_gpr_4,
  output [31:0] io_commit_gpr_5,
  output [31:0] io_commit_gpr_6,
  output [31:0] io_commit_gpr_7,
  output [31:0] io_commit_gpr_8,
  output [31:0] io_commit_gpr_9,
  output [31:0] io_commit_gpr_10,
  output [31:0] io_commit_gpr_11,
  output [31:0] io_commit_gpr_12,
  output [31:0] io_commit_gpr_13,
  output [31:0] io_commit_gpr_14,
  output [31:0] io_commit_gpr_15,
  output [31:0] io_commit_gpr_16,
  output [31:0] io_commit_gpr_17,
  output [31:0] io_commit_gpr_18,
  output [31:0] io_commit_gpr_19,
  output [31:0] io_commit_gpr_20,
  output [31:0] io_commit_gpr_21,
  output [31:0] io_commit_gpr_22,
  output [31:0] io_commit_gpr_23,
  output [31:0] io_commit_gpr_24,
  output [31:0] io_commit_gpr_25,
  output [31:0] io_commit_gpr_26,
  output [31:0] io_commit_gpr_27,
  output [31:0] io_commit_gpr_28,
  output [31:0] io_commit_gpr_29,
  output [31:0] io_commit_gpr_30,
  output [31:0] io_commit_gpr_31,
  output [4:0]  io_commit_rd_idx,
  output [31:0] io_commit_wdata,
  output        io_commit_wen,
  input         io_ex_flush_valid
);
  reg [7:0] wbids [0:31]; // @[rf.scala 21:18]
  reg [31:0] _RAND_0;
  wire [7:0] wbids__T_183_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_183_addr; // @[rf.scala 21:18]
  wire [7:0] wbids__T_1_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_1_addr; // @[rf.scala 21:18]
  wire  wbids__T_1_mask; // @[rf.scala 21:18]
  wire  wbids__T_1_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_5_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_5_addr; // @[rf.scala 21:18]
  wire  wbids__T_5_mask; // @[rf.scala 21:18]
  wire  wbids__T_5_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_9_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_9_addr; // @[rf.scala 21:18]
  wire  wbids__T_9_mask; // @[rf.scala 21:18]
  wire  wbids__T_9_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_13_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_13_addr; // @[rf.scala 21:18]
  wire  wbids__T_13_mask; // @[rf.scala 21:18]
  wire  wbids__T_13_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_17_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_17_addr; // @[rf.scala 21:18]
  wire  wbids__T_17_mask; // @[rf.scala 21:18]
  wire  wbids__T_17_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_21_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_21_addr; // @[rf.scala 21:18]
  wire  wbids__T_21_mask; // @[rf.scala 21:18]
  wire  wbids__T_21_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_25_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_25_addr; // @[rf.scala 21:18]
  wire  wbids__T_25_mask; // @[rf.scala 21:18]
  wire  wbids__T_25_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_29_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_29_addr; // @[rf.scala 21:18]
  wire  wbids__T_29_mask; // @[rf.scala 21:18]
  wire  wbids__T_29_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_33_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_33_addr; // @[rf.scala 21:18]
  wire  wbids__T_33_mask; // @[rf.scala 21:18]
  wire  wbids__T_33_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_37_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_37_addr; // @[rf.scala 21:18]
  wire  wbids__T_37_mask; // @[rf.scala 21:18]
  wire  wbids__T_37_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_41_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_41_addr; // @[rf.scala 21:18]
  wire  wbids__T_41_mask; // @[rf.scala 21:18]
  wire  wbids__T_41_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_45_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_45_addr; // @[rf.scala 21:18]
  wire  wbids__T_45_mask; // @[rf.scala 21:18]
  wire  wbids__T_45_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_49_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_49_addr; // @[rf.scala 21:18]
  wire  wbids__T_49_mask; // @[rf.scala 21:18]
  wire  wbids__T_49_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_53_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_53_addr; // @[rf.scala 21:18]
  wire  wbids__T_53_mask; // @[rf.scala 21:18]
  wire  wbids__T_53_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_57_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_57_addr; // @[rf.scala 21:18]
  wire  wbids__T_57_mask; // @[rf.scala 21:18]
  wire  wbids__T_57_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_61_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_61_addr; // @[rf.scala 21:18]
  wire  wbids__T_61_mask; // @[rf.scala 21:18]
  wire  wbids__T_61_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_65_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_65_addr; // @[rf.scala 21:18]
  wire  wbids__T_65_mask; // @[rf.scala 21:18]
  wire  wbids__T_65_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_69_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_69_addr; // @[rf.scala 21:18]
  wire  wbids__T_69_mask; // @[rf.scala 21:18]
  wire  wbids__T_69_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_73_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_73_addr; // @[rf.scala 21:18]
  wire  wbids__T_73_mask; // @[rf.scala 21:18]
  wire  wbids__T_73_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_77_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_77_addr; // @[rf.scala 21:18]
  wire  wbids__T_77_mask; // @[rf.scala 21:18]
  wire  wbids__T_77_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_81_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_81_addr; // @[rf.scala 21:18]
  wire  wbids__T_81_mask; // @[rf.scala 21:18]
  wire  wbids__T_81_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_85_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_85_addr; // @[rf.scala 21:18]
  wire  wbids__T_85_mask; // @[rf.scala 21:18]
  wire  wbids__T_85_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_89_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_89_addr; // @[rf.scala 21:18]
  wire  wbids__T_89_mask; // @[rf.scala 21:18]
  wire  wbids__T_89_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_93_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_93_addr; // @[rf.scala 21:18]
  wire  wbids__T_93_mask; // @[rf.scala 21:18]
  wire  wbids__T_93_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_97_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_97_addr; // @[rf.scala 21:18]
  wire  wbids__T_97_mask; // @[rf.scala 21:18]
  wire  wbids__T_97_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_101_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_101_addr; // @[rf.scala 21:18]
  wire  wbids__T_101_mask; // @[rf.scala 21:18]
  wire  wbids__T_101_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_105_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_105_addr; // @[rf.scala 21:18]
  wire  wbids__T_105_mask; // @[rf.scala 21:18]
  wire  wbids__T_105_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_109_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_109_addr; // @[rf.scala 21:18]
  wire  wbids__T_109_mask; // @[rf.scala 21:18]
  wire  wbids__T_109_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_113_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_113_addr; // @[rf.scala 21:18]
  wire  wbids__T_113_mask; // @[rf.scala 21:18]
  wire  wbids__T_113_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_117_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_117_addr; // @[rf.scala 21:18]
  wire  wbids__T_117_mask; // @[rf.scala 21:18]
  wire  wbids__T_117_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_121_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_121_addr; // @[rf.scala 21:18]
  wire  wbids__T_121_mask; // @[rf.scala 21:18]
  wire  wbids__T_121_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_125_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_125_addr; // @[rf.scala 21:18]
  wire  wbids__T_125_mask; // @[rf.scala 21:18]
  wire  wbids__T_125_en; // @[rf.scala 21:18]
  wire [7:0] wbids__T_194_data; // @[rf.scala 21:18]
  wire [4:0] wbids__T_194_addr; // @[rf.scala 21:18]
  wire  wbids__T_194_mask; // @[rf.scala 21:18]
  wire  wbids__T_194_en; // @[rf.scala 21:18]
  reg [31:0] wb_rf [0:31]; // @[rf.scala 22:18]
  reg [31:0] _RAND_1;
  wire [31:0] wb_rf__T_143_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_143_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_168_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_168_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_268_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_268_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_273_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_273_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_278_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_278_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_283_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_283_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_288_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_288_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_293_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_293_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_298_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_298_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_303_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_303_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_308_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_308_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_313_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_313_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_318_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_318_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_323_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_323_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_328_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_328_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_333_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_333_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_338_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_338_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_343_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_343_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_348_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_348_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_353_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_353_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_358_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_358_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_363_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_363_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_368_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_368_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_373_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_373_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_378_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_378_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_383_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_383_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_388_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_388_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_393_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_393_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_398_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_398_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_403_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_403_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_408_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_408_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_413_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_413_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_418_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_418_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_423_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_423_addr; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_4_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_4_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_4_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_4_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_8_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_8_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_8_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_8_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_12_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_12_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_12_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_12_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_16_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_16_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_16_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_16_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_20_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_20_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_20_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_20_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_24_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_24_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_24_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_24_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_28_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_28_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_28_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_28_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_32_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_32_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_32_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_32_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_36_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_36_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_36_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_36_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_40_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_40_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_40_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_40_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_44_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_44_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_44_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_44_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_48_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_48_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_48_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_48_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_52_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_52_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_52_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_52_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_56_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_56_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_56_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_56_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_60_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_60_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_60_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_60_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_64_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_64_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_64_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_64_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_68_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_68_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_68_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_68_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_72_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_72_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_72_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_72_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_76_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_76_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_76_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_76_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_80_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_80_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_80_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_80_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_84_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_84_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_84_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_84_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_88_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_88_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_88_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_88_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_92_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_92_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_92_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_92_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_96_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_96_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_96_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_96_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_100_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_100_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_100_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_100_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_104_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_104_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_104_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_104_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_108_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_108_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_108_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_108_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_112_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_112_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_112_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_112_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_116_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_116_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_116_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_116_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_120_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_120_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_120_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_120_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_124_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_124_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_124_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_124_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_128_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_128_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_128_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_128_en; // @[rf.scala 22:18]
  wire [31:0] wb_rf__T_182_data; // @[rf.scala 22:18]
  wire [4:0] wb_rf__T_182_addr; // @[rf.scala 22:18]
  wire  wb_rf__T_182_mask; // @[rf.scala 22:18]
  wire  wb_rf__T_182_en; // @[rf.scala 22:18]
  reg [31:0] bp_rf [0:31]; // @[rf.scala 23:18]
  reg [31:0] _RAND_2;
  wire [31:0] bp_rf__T_149_data; // @[rf.scala 23:18]
  wire [4:0] bp_rf__T_149_addr; // @[rf.scala 23:18]
  wire [31:0] bp_rf__T_174_data; // @[rf.scala 23:18]
  wire [4:0] bp_rf__T_174_addr; // @[rf.scala 23:18]
  wire [31:0] bp_rf__T_190_data; // @[rf.scala 23:18]
  wire [4:0] bp_rf__T_190_addr; // @[rf.scala 23:18]
  wire  bp_rf__T_190_mask; // @[rf.scala 23:18]
  wire  bp_rf__T_190_en; // @[rf.scala 23:18]
  reg  rf_dirtys [0:31]; // @[rf.scala 24:22]
  reg [31:0] _RAND_3;
  wire  rf_dirtys__T_129_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_129_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_141_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_141_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_154_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_154_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_166_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_166_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_2_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_2_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_2_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_2_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_6_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_6_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_6_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_6_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_10_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_10_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_10_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_10_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_14_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_14_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_14_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_14_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_18_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_18_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_18_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_18_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_22_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_22_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_22_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_22_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_26_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_26_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_26_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_26_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_30_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_30_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_30_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_30_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_34_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_34_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_34_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_34_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_38_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_38_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_38_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_38_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_42_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_42_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_42_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_42_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_46_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_46_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_46_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_46_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_50_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_50_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_50_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_50_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_54_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_54_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_54_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_54_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_58_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_58_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_58_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_58_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_62_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_62_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_62_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_62_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_66_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_66_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_66_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_66_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_70_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_70_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_70_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_70_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_74_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_74_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_74_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_74_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_78_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_78_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_78_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_78_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_82_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_82_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_82_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_82_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_86_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_86_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_86_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_86_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_90_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_90_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_90_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_90_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_94_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_94_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_94_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_94_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_98_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_98_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_98_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_98_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_102_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_102_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_102_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_102_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_106_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_106_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_106_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_106_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_110_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_110_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_110_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_110_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_114_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_114_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_114_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_114_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_118_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_118_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_118_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_118_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_122_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_122_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_122_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_122_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_126_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_126_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_126_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_126_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_185_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_185_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_185_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_185_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_192_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_192_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_192_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_192_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_195_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_195_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_195_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_195_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_197_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_197_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_197_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_197_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_199_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_199_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_199_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_199_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_201_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_201_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_201_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_201_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_203_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_203_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_203_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_203_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_205_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_205_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_205_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_205_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_207_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_207_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_207_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_207_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_209_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_209_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_209_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_209_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_211_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_211_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_211_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_211_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_213_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_213_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_213_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_213_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_215_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_215_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_215_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_215_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_217_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_217_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_217_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_217_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_219_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_219_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_219_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_219_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_221_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_221_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_221_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_221_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_223_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_223_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_223_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_223_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_225_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_225_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_225_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_225_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_227_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_227_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_227_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_227_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_229_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_229_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_229_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_229_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_231_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_231_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_231_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_231_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_233_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_233_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_233_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_233_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_235_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_235_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_235_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_235_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_237_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_237_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_237_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_237_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_239_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_239_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_239_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_239_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_241_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_241_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_241_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_241_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_243_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_243_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_243_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_243_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_245_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_245_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_245_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_245_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_247_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_247_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_247_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_247_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_249_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_249_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_249_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_249_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_251_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_251_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_251_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_251_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_253_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_253_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_253_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_253_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_255_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_255_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_255_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_255_en; // @[rf.scala 24:22]
  wire  rf_dirtys__T_257_data; // @[rf.scala 24:22]
  wire [4:0] rf_dirtys__T_257_addr; // @[rf.scala 24:22]
  wire  rf_dirtys__T_257_mask; // @[rf.scala 24:22]
  wire  rf_dirtys__T_257_en; // @[rf.scala 24:22]
  reg  bp_readys [0:31]; // @[rf.scala 25:22]
  reg [31:0] _RAND_4;
  wire  bp_readys__T_131_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_131_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_148_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_148_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_156_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_156_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_173_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_173_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_3_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_3_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_3_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_3_en; // @[rf.scala 25:22]
  wire  bp_readys__T_7_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_7_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_7_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_7_en; // @[rf.scala 25:22]
  wire  bp_readys__T_11_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_11_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_11_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_11_en; // @[rf.scala 25:22]
  wire  bp_readys__T_15_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_15_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_15_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_15_en; // @[rf.scala 25:22]
  wire  bp_readys__T_19_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_19_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_19_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_19_en; // @[rf.scala 25:22]
  wire  bp_readys__T_23_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_23_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_23_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_23_en; // @[rf.scala 25:22]
  wire  bp_readys__T_27_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_27_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_27_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_27_en; // @[rf.scala 25:22]
  wire  bp_readys__T_31_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_31_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_31_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_31_en; // @[rf.scala 25:22]
  wire  bp_readys__T_35_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_35_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_35_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_35_en; // @[rf.scala 25:22]
  wire  bp_readys__T_39_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_39_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_39_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_39_en; // @[rf.scala 25:22]
  wire  bp_readys__T_43_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_43_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_43_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_43_en; // @[rf.scala 25:22]
  wire  bp_readys__T_47_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_47_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_47_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_47_en; // @[rf.scala 25:22]
  wire  bp_readys__T_51_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_51_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_51_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_51_en; // @[rf.scala 25:22]
  wire  bp_readys__T_55_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_55_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_55_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_55_en; // @[rf.scala 25:22]
  wire  bp_readys__T_59_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_59_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_59_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_59_en; // @[rf.scala 25:22]
  wire  bp_readys__T_63_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_63_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_63_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_63_en; // @[rf.scala 25:22]
  wire  bp_readys__T_67_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_67_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_67_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_67_en; // @[rf.scala 25:22]
  wire  bp_readys__T_71_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_71_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_71_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_71_en; // @[rf.scala 25:22]
  wire  bp_readys__T_75_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_75_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_75_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_75_en; // @[rf.scala 25:22]
  wire  bp_readys__T_79_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_79_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_79_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_79_en; // @[rf.scala 25:22]
  wire  bp_readys__T_83_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_83_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_83_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_83_en; // @[rf.scala 25:22]
  wire  bp_readys__T_87_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_87_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_87_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_87_en; // @[rf.scala 25:22]
  wire  bp_readys__T_91_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_91_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_91_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_91_en; // @[rf.scala 25:22]
  wire  bp_readys__T_95_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_95_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_95_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_95_en; // @[rf.scala 25:22]
  wire  bp_readys__T_99_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_99_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_99_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_99_en; // @[rf.scala 25:22]
  wire  bp_readys__T_103_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_103_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_103_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_103_en; // @[rf.scala 25:22]
  wire  bp_readys__T_107_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_107_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_107_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_107_en; // @[rf.scala 25:22]
  wire  bp_readys__T_111_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_111_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_111_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_111_en; // @[rf.scala 25:22]
  wire  bp_readys__T_115_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_115_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_115_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_115_en; // @[rf.scala 25:22]
  wire  bp_readys__T_119_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_119_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_119_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_119_en; // @[rf.scala 25:22]
  wire  bp_readys__T_123_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_123_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_123_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_123_en; // @[rf.scala 25:22]
  wire  bp_readys__T_127_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_127_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_127_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_127_en; // @[rf.scala 25:22]
  wire  bp_readys__T_191_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_191_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_191_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_191_en; // @[rf.scala 25:22]
  wire  bp_readys__T_193_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_193_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_193_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_193_en; // @[rf.scala 25:22]
  wire  bp_readys__T_196_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_196_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_196_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_196_en; // @[rf.scala 25:22]
  wire  bp_readys__T_198_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_198_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_198_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_198_en; // @[rf.scala 25:22]
  wire  bp_readys__T_200_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_200_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_200_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_200_en; // @[rf.scala 25:22]
  wire  bp_readys__T_202_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_202_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_202_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_202_en; // @[rf.scala 25:22]
  wire  bp_readys__T_204_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_204_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_204_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_204_en; // @[rf.scala 25:22]
  wire  bp_readys__T_206_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_206_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_206_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_206_en; // @[rf.scala 25:22]
  wire  bp_readys__T_208_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_208_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_208_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_208_en; // @[rf.scala 25:22]
  wire  bp_readys__T_210_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_210_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_210_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_210_en; // @[rf.scala 25:22]
  wire  bp_readys__T_212_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_212_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_212_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_212_en; // @[rf.scala 25:22]
  wire  bp_readys__T_214_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_214_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_214_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_214_en; // @[rf.scala 25:22]
  wire  bp_readys__T_216_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_216_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_216_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_216_en; // @[rf.scala 25:22]
  wire  bp_readys__T_218_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_218_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_218_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_218_en; // @[rf.scala 25:22]
  wire  bp_readys__T_220_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_220_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_220_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_220_en; // @[rf.scala 25:22]
  wire  bp_readys__T_222_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_222_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_222_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_222_en; // @[rf.scala 25:22]
  wire  bp_readys__T_224_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_224_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_224_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_224_en; // @[rf.scala 25:22]
  wire  bp_readys__T_226_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_226_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_226_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_226_en; // @[rf.scala 25:22]
  wire  bp_readys__T_228_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_228_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_228_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_228_en; // @[rf.scala 25:22]
  wire  bp_readys__T_230_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_230_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_230_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_230_en; // @[rf.scala 25:22]
  wire  bp_readys__T_232_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_232_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_232_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_232_en; // @[rf.scala 25:22]
  wire  bp_readys__T_234_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_234_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_234_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_234_en; // @[rf.scala 25:22]
  wire  bp_readys__T_236_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_236_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_236_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_236_en; // @[rf.scala 25:22]
  wire  bp_readys__T_238_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_238_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_238_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_238_en; // @[rf.scala 25:22]
  wire  bp_readys__T_240_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_240_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_240_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_240_en; // @[rf.scala 25:22]
  wire  bp_readys__T_242_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_242_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_242_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_242_en; // @[rf.scala 25:22]
  wire  bp_readys__T_244_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_244_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_244_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_244_en; // @[rf.scala 25:22]
  wire  bp_readys__T_246_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_246_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_246_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_246_en; // @[rf.scala 25:22]
  wire  bp_readys__T_248_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_248_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_248_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_248_en; // @[rf.scala 25:22]
  wire  bp_readys__T_250_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_250_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_250_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_250_en; // @[rf.scala 25:22]
  wire  bp_readys__T_252_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_252_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_252_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_252_en; // @[rf.scala 25:22]
  wire  bp_readys__T_254_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_254_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_254_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_254_en; // @[rf.scala 25:22]
  wire  bp_readys__T_256_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_256_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_256_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_256_en; // @[rf.scala 25:22]
  wire  bp_readys__T_258_data; // @[rf.scala 25:22]
  wire [4:0] bp_readys__T_258_addr; // @[rf.scala 25:22]
  wire  bp_readys__T_258_mask; // @[rf.scala 25:22]
  wire  bp_readys__T_258_en; // @[rf.scala 25:22]
  wire  _T_130 = ~rf_dirtys__T_129_data; // @[rf.scala 37:33]
  wire  _T_132 = _T_130 | bp_readys__T_131_data; // @[rf.scala 37:49]
  wire  _T_133 = io_bp_valid & io_bp_bits_v; // @[rf.scala 36:44]
  wire  _T_134 = _T_133 & io_bp_bits_wen; // @[rf.scala 36:60]
  wire  _T_135 = io_bp_bits_rd_idx == io_rfio_rs_idx; // @[rf.scala 36:99]
  wire  _T_136 = _T_134 & _T_135; // @[rf.scala 36:78]
  wire  _T_137 = _T_132 | _T_136; // @[rf.scala 37:67]
  wire  _T_138 = io_rfio_rs_idx == 5'h0; // @[rf.scala 37:95]
  wire  _T_142 = ~rf_dirtys__T_141_data; // @[rf.scala 40:5]
  wire [31:0] _T_150 = bp_readys__T_148_data ? bp_rf__T_149_data : 32'h0; // @[Mux.scala 87:16]
  wire [31:0] _T_151 = _T_136 ? io_bp_bits_data : _T_150; // @[Mux.scala 87:16]
  wire [31:0] _T_152 = _T_142 ? wb_rf__T_143_data : _T_151; // @[Mux.scala 87:16]
  wire  _T_155 = ~rf_dirtys__T_154_data; // @[rf.scala 37:33]
  wire  _T_157 = _T_155 | bp_readys__T_156_data; // @[rf.scala 37:49]
  wire  _T_160 = io_bp_bits_rd_idx == io_rfio_rt_idx; // @[rf.scala 36:99]
  wire  _T_161 = _T_134 & _T_160; // @[rf.scala 36:78]
  wire  _T_162 = _T_157 | _T_161; // @[rf.scala 37:67]
  wire  _T_163 = io_rfio_rt_idx == 5'h0; // @[rf.scala 37:95]
  wire  _T_167 = ~rf_dirtys__T_166_data; // @[rf.scala 40:5]
  wire [31:0] _T_175 = bp_readys__T_173_data ? bp_rf__T_174_data : 32'h0; // @[Mux.scala 87:16]
  wire [31:0] _T_176 = _T_161 ? io_bp_bits_data : _T_175; // @[Mux.scala 87:16]
  wire [31:0] _T_177 = _T_167 ? wb_rf__T_168_data : _T_176; // @[Mux.scala 87:16]
  wire  _T_179 = io_wb_valid & io_wb_bits_v; // @[rf.scala 50:21]
  wire  _T_180 = io_wb_bits_rd_idx != 5'h0; // @[rf.scala 51:47]
  wire  _T_181 = io_wb_bits_wen & _T_180; // @[rf.scala 51:26]
  wire  _T_184 = wbids__T_183_data == io_wb_bits_id; // @[rf.scala 54:36]
  wire  _T_188 = io_bp_bits_rd_idx != 5'h0; // @[rf.scala 60:23]
  wire [15:0] _T_260 = {io_wb_bits_instr_rd_idx,io_wb_bits_instr_shamt,io_wb_bits_instr_func}; // @[rf.scala 81:39]
  wire [15:0] _T_262 = {io_wb_bits_instr_op,io_wb_bits_instr_rs_idx,io_wb_bits_instr_rt_idx}; // @[rf.scala 81:39]
  wire  _T_265 = io_wb_valid & io_wb_bits_wen; // @[rf.scala 87:41]
  wire  _T_266 = io_wb_bits_rd_idx == 5'h0; // @[rf.scala 87:80]
  wire  _T_267 = _T_265 & _T_266; // @[rf.scala 87:59]
  wire  _T_271 = io_wb_bits_rd_idx == 5'h1; // @[rf.scala 87:80]
  wire  _T_272 = _T_265 & _T_271; // @[rf.scala 87:59]
  wire  _T_276 = io_wb_bits_rd_idx == 5'h2; // @[rf.scala 87:80]
  wire  _T_277 = _T_265 & _T_276; // @[rf.scala 87:59]
  wire  _T_281 = io_wb_bits_rd_idx == 5'h3; // @[rf.scala 87:80]
  wire  _T_282 = _T_265 & _T_281; // @[rf.scala 87:59]
  wire  _T_286 = io_wb_bits_rd_idx == 5'h4; // @[rf.scala 87:80]
  wire  _T_287 = _T_265 & _T_286; // @[rf.scala 87:59]
  wire  _T_291 = io_wb_bits_rd_idx == 5'h5; // @[rf.scala 87:80]
  wire  _T_292 = _T_265 & _T_291; // @[rf.scala 87:59]
  wire  _T_296 = io_wb_bits_rd_idx == 5'h6; // @[rf.scala 87:80]
  wire  _T_297 = _T_265 & _T_296; // @[rf.scala 87:59]
  wire  _T_301 = io_wb_bits_rd_idx == 5'h7; // @[rf.scala 87:80]
  wire  _T_302 = _T_265 & _T_301; // @[rf.scala 87:59]
  wire  _T_306 = io_wb_bits_rd_idx == 5'h8; // @[rf.scala 87:80]
  wire  _T_307 = _T_265 & _T_306; // @[rf.scala 87:59]
  wire  _T_311 = io_wb_bits_rd_idx == 5'h9; // @[rf.scala 87:80]
  wire  _T_312 = _T_265 & _T_311; // @[rf.scala 87:59]
  wire  _T_316 = io_wb_bits_rd_idx == 5'ha; // @[rf.scala 87:80]
  wire  _T_317 = _T_265 & _T_316; // @[rf.scala 87:59]
  wire  _T_321 = io_wb_bits_rd_idx == 5'hb; // @[rf.scala 87:80]
  wire  _T_322 = _T_265 & _T_321; // @[rf.scala 87:59]
  wire  _T_326 = io_wb_bits_rd_idx == 5'hc; // @[rf.scala 87:80]
  wire  _T_327 = _T_265 & _T_326; // @[rf.scala 87:59]
  wire  _T_331 = io_wb_bits_rd_idx == 5'hd; // @[rf.scala 87:80]
  wire  _T_332 = _T_265 & _T_331; // @[rf.scala 87:59]
  wire  _T_336 = io_wb_bits_rd_idx == 5'he; // @[rf.scala 87:80]
  wire  _T_337 = _T_265 & _T_336; // @[rf.scala 87:59]
  wire  _T_341 = io_wb_bits_rd_idx == 5'hf; // @[rf.scala 87:80]
  wire  _T_342 = _T_265 & _T_341; // @[rf.scala 87:59]
  wire  _T_346 = io_wb_bits_rd_idx == 5'h10; // @[rf.scala 87:80]
  wire  _T_347 = _T_265 & _T_346; // @[rf.scala 87:59]
  wire  _T_351 = io_wb_bits_rd_idx == 5'h11; // @[rf.scala 87:80]
  wire  _T_352 = _T_265 & _T_351; // @[rf.scala 87:59]
  wire  _T_356 = io_wb_bits_rd_idx == 5'h12; // @[rf.scala 87:80]
  wire  _T_357 = _T_265 & _T_356; // @[rf.scala 87:59]
  wire  _T_361 = io_wb_bits_rd_idx == 5'h13; // @[rf.scala 87:80]
  wire  _T_362 = _T_265 & _T_361; // @[rf.scala 87:59]
  wire  _T_366 = io_wb_bits_rd_idx == 5'h14; // @[rf.scala 87:80]
  wire  _T_367 = _T_265 & _T_366; // @[rf.scala 87:59]
  wire  _T_371 = io_wb_bits_rd_idx == 5'h15; // @[rf.scala 87:80]
  wire  _T_372 = _T_265 & _T_371; // @[rf.scala 87:59]
  wire  _T_376 = io_wb_bits_rd_idx == 5'h16; // @[rf.scala 87:80]
  wire  _T_377 = _T_265 & _T_376; // @[rf.scala 87:59]
  wire  _T_381 = io_wb_bits_rd_idx == 5'h17; // @[rf.scala 87:80]
  wire  _T_382 = _T_265 & _T_381; // @[rf.scala 87:59]
  wire  _T_386 = io_wb_bits_rd_idx == 5'h18; // @[rf.scala 87:80]
  wire  _T_387 = _T_265 & _T_386; // @[rf.scala 87:59]
  wire  _T_391 = io_wb_bits_rd_idx == 5'h19; // @[rf.scala 87:80]
  wire  _T_392 = _T_265 & _T_391; // @[rf.scala 87:59]
  wire  _T_396 = io_wb_bits_rd_idx == 5'h1a; // @[rf.scala 87:80]
  wire  _T_397 = _T_265 & _T_396; // @[rf.scala 87:59]
  wire  _T_401 = io_wb_bits_rd_idx == 5'h1b; // @[rf.scala 87:80]
  wire  _T_402 = _T_265 & _T_401; // @[rf.scala 87:59]
  wire  _T_406 = io_wb_bits_rd_idx == 5'h1c; // @[rf.scala 87:80]
  wire  _T_407 = _T_265 & _T_406; // @[rf.scala 87:59]
  wire  _T_411 = io_wb_bits_rd_idx == 5'h1d; // @[rf.scala 87:80]
  wire  _T_412 = _T_265 & _T_411; // @[rf.scala 87:59]
  wire  _T_416 = io_wb_bits_rd_idx == 5'h1e; // @[rf.scala 87:80]
  wire  _T_417 = _T_265 & _T_416; // @[rf.scala 87:59]
  wire  _T_421 = io_wb_bits_rd_idx == 5'h1f; // @[rf.scala 87:80]
  wire  _T_422 = _T_265 & _T_421; // @[rf.scala 87:59]
  assign wbids__T_183_addr = io_wb_bits_rd_idx;
  assign wbids__T_183_data = wbids[wbids__T_183_addr]; // @[rf.scala 21:18]
  assign wbids__T_1_data = 8'h0;
  assign wbids__T_1_addr = 5'h0;
  assign wbids__T_1_mask = 1'h1;
  assign wbids__T_1_en = reset;
  assign wbids__T_5_data = 8'h0;
  assign wbids__T_5_addr = 5'h1;
  assign wbids__T_5_mask = 1'h1;
  assign wbids__T_5_en = reset;
  assign wbids__T_9_data = 8'h0;
  assign wbids__T_9_addr = 5'h2;
  assign wbids__T_9_mask = 1'h1;
  assign wbids__T_9_en = reset;
  assign wbids__T_13_data = 8'h0;
  assign wbids__T_13_addr = 5'h3;
  assign wbids__T_13_mask = 1'h1;
  assign wbids__T_13_en = reset;
  assign wbids__T_17_data = 8'h0;
  assign wbids__T_17_addr = 5'h4;
  assign wbids__T_17_mask = 1'h1;
  assign wbids__T_17_en = reset;
  assign wbids__T_21_data = 8'h0;
  assign wbids__T_21_addr = 5'h5;
  assign wbids__T_21_mask = 1'h1;
  assign wbids__T_21_en = reset;
  assign wbids__T_25_data = 8'h0;
  assign wbids__T_25_addr = 5'h6;
  assign wbids__T_25_mask = 1'h1;
  assign wbids__T_25_en = reset;
  assign wbids__T_29_data = 8'h0;
  assign wbids__T_29_addr = 5'h7;
  assign wbids__T_29_mask = 1'h1;
  assign wbids__T_29_en = reset;
  assign wbids__T_33_data = 8'h0;
  assign wbids__T_33_addr = 5'h8;
  assign wbids__T_33_mask = 1'h1;
  assign wbids__T_33_en = reset;
  assign wbids__T_37_data = 8'h0;
  assign wbids__T_37_addr = 5'h9;
  assign wbids__T_37_mask = 1'h1;
  assign wbids__T_37_en = reset;
  assign wbids__T_41_data = 8'h0;
  assign wbids__T_41_addr = 5'ha;
  assign wbids__T_41_mask = 1'h1;
  assign wbids__T_41_en = reset;
  assign wbids__T_45_data = 8'h0;
  assign wbids__T_45_addr = 5'hb;
  assign wbids__T_45_mask = 1'h1;
  assign wbids__T_45_en = reset;
  assign wbids__T_49_data = 8'h0;
  assign wbids__T_49_addr = 5'hc;
  assign wbids__T_49_mask = 1'h1;
  assign wbids__T_49_en = reset;
  assign wbids__T_53_data = 8'h0;
  assign wbids__T_53_addr = 5'hd;
  assign wbids__T_53_mask = 1'h1;
  assign wbids__T_53_en = reset;
  assign wbids__T_57_data = 8'h0;
  assign wbids__T_57_addr = 5'he;
  assign wbids__T_57_mask = 1'h1;
  assign wbids__T_57_en = reset;
  assign wbids__T_61_data = 8'h0;
  assign wbids__T_61_addr = 5'hf;
  assign wbids__T_61_mask = 1'h1;
  assign wbids__T_61_en = reset;
  assign wbids__T_65_data = 8'h0;
  assign wbids__T_65_addr = 5'h10;
  assign wbids__T_65_mask = 1'h1;
  assign wbids__T_65_en = reset;
  assign wbids__T_69_data = 8'h0;
  assign wbids__T_69_addr = 5'h11;
  assign wbids__T_69_mask = 1'h1;
  assign wbids__T_69_en = reset;
  assign wbids__T_73_data = 8'h0;
  assign wbids__T_73_addr = 5'h12;
  assign wbids__T_73_mask = 1'h1;
  assign wbids__T_73_en = reset;
  assign wbids__T_77_data = 8'h0;
  assign wbids__T_77_addr = 5'h13;
  assign wbids__T_77_mask = 1'h1;
  assign wbids__T_77_en = reset;
  assign wbids__T_81_data = 8'h0;
  assign wbids__T_81_addr = 5'h14;
  assign wbids__T_81_mask = 1'h1;
  assign wbids__T_81_en = reset;
  assign wbids__T_85_data = 8'h0;
  assign wbids__T_85_addr = 5'h15;
  assign wbids__T_85_mask = 1'h1;
  assign wbids__T_85_en = reset;
  assign wbids__T_89_data = 8'h0;
  assign wbids__T_89_addr = 5'h16;
  assign wbids__T_89_mask = 1'h1;
  assign wbids__T_89_en = reset;
  assign wbids__T_93_data = 8'h0;
  assign wbids__T_93_addr = 5'h17;
  assign wbids__T_93_mask = 1'h1;
  assign wbids__T_93_en = reset;
  assign wbids__T_97_data = 8'h0;
  assign wbids__T_97_addr = 5'h18;
  assign wbids__T_97_mask = 1'h1;
  assign wbids__T_97_en = reset;
  assign wbids__T_101_data = 8'h0;
  assign wbids__T_101_addr = 5'h19;
  assign wbids__T_101_mask = 1'h1;
  assign wbids__T_101_en = reset;
  assign wbids__T_105_data = 8'h0;
  assign wbids__T_105_addr = 5'h1a;
  assign wbids__T_105_mask = 1'h1;
  assign wbids__T_105_en = reset;
  assign wbids__T_109_data = 8'h0;
  assign wbids__T_109_addr = 5'h1b;
  assign wbids__T_109_mask = 1'h1;
  assign wbids__T_109_en = reset;
  assign wbids__T_113_data = 8'h0;
  assign wbids__T_113_addr = 5'h1c;
  assign wbids__T_113_mask = 1'h1;
  assign wbids__T_113_en = reset;
  assign wbids__T_117_data = 8'h0;
  assign wbids__T_117_addr = 5'h1d;
  assign wbids__T_117_mask = 1'h1;
  assign wbids__T_117_en = reset;
  assign wbids__T_121_data = 8'h0;
  assign wbids__T_121_addr = 5'h1e;
  assign wbids__T_121_mask = 1'h1;
  assign wbids__T_121_en = reset;
  assign wbids__T_125_data = 8'h0;
  assign wbids__T_125_addr = 5'h1f;
  assign wbids__T_125_mask = 1'h1;
  assign wbids__T_125_en = reset;
  assign wbids__T_194_data = io_rfio_wid;
  assign wbids__T_194_addr = io_rfio_rd_idx;
  assign wbids__T_194_mask = 1'h1;
  assign wbids__T_194_en = io_rfio_wen;
  assign wb_rf__T_143_addr = io_rfio_rs_idx;
  assign wb_rf__T_143_data = wb_rf[wb_rf__T_143_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_168_addr = io_rfio_rt_idx;
  assign wb_rf__T_168_data = wb_rf[wb_rf__T_168_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_268_addr = 5'h0;
  assign wb_rf__T_268_data = wb_rf[wb_rf__T_268_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_273_addr = 5'h1;
  assign wb_rf__T_273_data = wb_rf[wb_rf__T_273_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_278_addr = 5'h2;
  assign wb_rf__T_278_data = wb_rf[wb_rf__T_278_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_283_addr = 5'h3;
  assign wb_rf__T_283_data = wb_rf[wb_rf__T_283_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_288_addr = 5'h4;
  assign wb_rf__T_288_data = wb_rf[wb_rf__T_288_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_293_addr = 5'h5;
  assign wb_rf__T_293_data = wb_rf[wb_rf__T_293_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_298_addr = 5'h6;
  assign wb_rf__T_298_data = wb_rf[wb_rf__T_298_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_303_addr = 5'h7;
  assign wb_rf__T_303_data = wb_rf[wb_rf__T_303_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_308_addr = 5'h8;
  assign wb_rf__T_308_data = wb_rf[wb_rf__T_308_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_313_addr = 5'h9;
  assign wb_rf__T_313_data = wb_rf[wb_rf__T_313_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_318_addr = 5'ha;
  assign wb_rf__T_318_data = wb_rf[wb_rf__T_318_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_323_addr = 5'hb;
  assign wb_rf__T_323_data = wb_rf[wb_rf__T_323_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_328_addr = 5'hc;
  assign wb_rf__T_328_data = wb_rf[wb_rf__T_328_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_333_addr = 5'hd;
  assign wb_rf__T_333_data = wb_rf[wb_rf__T_333_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_338_addr = 5'he;
  assign wb_rf__T_338_data = wb_rf[wb_rf__T_338_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_343_addr = 5'hf;
  assign wb_rf__T_343_data = wb_rf[wb_rf__T_343_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_348_addr = 5'h10;
  assign wb_rf__T_348_data = wb_rf[wb_rf__T_348_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_353_addr = 5'h11;
  assign wb_rf__T_353_data = wb_rf[wb_rf__T_353_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_358_addr = 5'h12;
  assign wb_rf__T_358_data = wb_rf[wb_rf__T_358_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_363_addr = 5'h13;
  assign wb_rf__T_363_data = wb_rf[wb_rf__T_363_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_368_addr = 5'h14;
  assign wb_rf__T_368_data = wb_rf[wb_rf__T_368_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_373_addr = 5'h15;
  assign wb_rf__T_373_data = wb_rf[wb_rf__T_373_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_378_addr = 5'h16;
  assign wb_rf__T_378_data = wb_rf[wb_rf__T_378_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_383_addr = 5'h17;
  assign wb_rf__T_383_data = wb_rf[wb_rf__T_383_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_388_addr = 5'h18;
  assign wb_rf__T_388_data = wb_rf[wb_rf__T_388_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_393_addr = 5'h19;
  assign wb_rf__T_393_data = wb_rf[wb_rf__T_393_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_398_addr = 5'h1a;
  assign wb_rf__T_398_data = wb_rf[wb_rf__T_398_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_403_addr = 5'h1b;
  assign wb_rf__T_403_data = wb_rf[wb_rf__T_403_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_408_addr = 5'h1c;
  assign wb_rf__T_408_data = wb_rf[wb_rf__T_408_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_413_addr = 5'h1d;
  assign wb_rf__T_413_data = wb_rf[wb_rf__T_413_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_418_addr = 5'h1e;
  assign wb_rf__T_418_data = wb_rf[wb_rf__T_418_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_423_addr = 5'h1f;
  assign wb_rf__T_423_data = wb_rf[wb_rf__T_423_addr]; // @[rf.scala 22:18]
  assign wb_rf__T_4_data = 32'h0;
  assign wb_rf__T_4_addr = 5'h0;
  assign wb_rf__T_4_mask = 1'h1;
  assign wb_rf__T_4_en = reset;
  assign wb_rf__T_8_data = 32'h0;
  assign wb_rf__T_8_addr = 5'h1;
  assign wb_rf__T_8_mask = 1'h1;
  assign wb_rf__T_8_en = reset;
  assign wb_rf__T_12_data = 32'h0;
  assign wb_rf__T_12_addr = 5'h2;
  assign wb_rf__T_12_mask = 1'h1;
  assign wb_rf__T_12_en = reset;
  assign wb_rf__T_16_data = 32'h0;
  assign wb_rf__T_16_addr = 5'h3;
  assign wb_rf__T_16_mask = 1'h1;
  assign wb_rf__T_16_en = reset;
  assign wb_rf__T_20_data = 32'h0;
  assign wb_rf__T_20_addr = 5'h4;
  assign wb_rf__T_20_mask = 1'h1;
  assign wb_rf__T_20_en = reset;
  assign wb_rf__T_24_data = 32'h0;
  assign wb_rf__T_24_addr = 5'h5;
  assign wb_rf__T_24_mask = 1'h1;
  assign wb_rf__T_24_en = reset;
  assign wb_rf__T_28_data = 32'h0;
  assign wb_rf__T_28_addr = 5'h6;
  assign wb_rf__T_28_mask = 1'h1;
  assign wb_rf__T_28_en = reset;
  assign wb_rf__T_32_data = 32'h0;
  assign wb_rf__T_32_addr = 5'h7;
  assign wb_rf__T_32_mask = 1'h1;
  assign wb_rf__T_32_en = reset;
  assign wb_rf__T_36_data = 32'h0;
  assign wb_rf__T_36_addr = 5'h8;
  assign wb_rf__T_36_mask = 1'h1;
  assign wb_rf__T_36_en = reset;
  assign wb_rf__T_40_data = 32'h0;
  assign wb_rf__T_40_addr = 5'h9;
  assign wb_rf__T_40_mask = 1'h1;
  assign wb_rf__T_40_en = reset;
  assign wb_rf__T_44_data = 32'h0;
  assign wb_rf__T_44_addr = 5'ha;
  assign wb_rf__T_44_mask = 1'h1;
  assign wb_rf__T_44_en = reset;
  assign wb_rf__T_48_data = 32'h0;
  assign wb_rf__T_48_addr = 5'hb;
  assign wb_rf__T_48_mask = 1'h1;
  assign wb_rf__T_48_en = reset;
  assign wb_rf__T_52_data = 32'h0;
  assign wb_rf__T_52_addr = 5'hc;
  assign wb_rf__T_52_mask = 1'h1;
  assign wb_rf__T_52_en = reset;
  assign wb_rf__T_56_data = 32'h0;
  assign wb_rf__T_56_addr = 5'hd;
  assign wb_rf__T_56_mask = 1'h1;
  assign wb_rf__T_56_en = reset;
  assign wb_rf__T_60_data = 32'h0;
  assign wb_rf__T_60_addr = 5'he;
  assign wb_rf__T_60_mask = 1'h1;
  assign wb_rf__T_60_en = reset;
  assign wb_rf__T_64_data = 32'h0;
  assign wb_rf__T_64_addr = 5'hf;
  assign wb_rf__T_64_mask = 1'h1;
  assign wb_rf__T_64_en = reset;
  assign wb_rf__T_68_data = 32'h0;
  assign wb_rf__T_68_addr = 5'h10;
  assign wb_rf__T_68_mask = 1'h1;
  assign wb_rf__T_68_en = reset;
  assign wb_rf__T_72_data = 32'h0;
  assign wb_rf__T_72_addr = 5'h11;
  assign wb_rf__T_72_mask = 1'h1;
  assign wb_rf__T_72_en = reset;
  assign wb_rf__T_76_data = 32'h0;
  assign wb_rf__T_76_addr = 5'h12;
  assign wb_rf__T_76_mask = 1'h1;
  assign wb_rf__T_76_en = reset;
  assign wb_rf__T_80_data = 32'h0;
  assign wb_rf__T_80_addr = 5'h13;
  assign wb_rf__T_80_mask = 1'h1;
  assign wb_rf__T_80_en = reset;
  assign wb_rf__T_84_data = 32'h0;
  assign wb_rf__T_84_addr = 5'h14;
  assign wb_rf__T_84_mask = 1'h1;
  assign wb_rf__T_84_en = reset;
  assign wb_rf__T_88_data = 32'h0;
  assign wb_rf__T_88_addr = 5'h15;
  assign wb_rf__T_88_mask = 1'h1;
  assign wb_rf__T_88_en = reset;
  assign wb_rf__T_92_data = 32'h0;
  assign wb_rf__T_92_addr = 5'h16;
  assign wb_rf__T_92_mask = 1'h1;
  assign wb_rf__T_92_en = reset;
  assign wb_rf__T_96_data = 32'h0;
  assign wb_rf__T_96_addr = 5'h17;
  assign wb_rf__T_96_mask = 1'h1;
  assign wb_rf__T_96_en = reset;
  assign wb_rf__T_100_data = 32'h0;
  assign wb_rf__T_100_addr = 5'h18;
  assign wb_rf__T_100_mask = 1'h1;
  assign wb_rf__T_100_en = reset;
  assign wb_rf__T_104_data = 32'h0;
  assign wb_rf__T_104_addr = 5'h19;
  assign wb_rf__T_104_mask = 1'h1;
  assign wb_rf__T_104_en = reset;
  assign wb_rf__T_108_data = 32'h0;
  assign wb_rf__T_108_addr = 5'h1a;
  assign wb_rf__T_108_mask = 1'h1;
  assign wb_rf__T_108_en = reset;
  assign wb_rf__T_112_data = 32'h0;
  assign wb_rf__T_112_addr = 5'h1b;
  assign wb_rf__T_112_mask = 1'h1;
  assign wb_rf__T_112_en = reset;
  assign wb_rf__T_116_data = 32'h0;
  assign wb_rf__T_116_addr = 5'h1c;
  assign wb_rf__T_116_mask = 1'h1;
  assign wb_rf__T_116_en = reset;
  assign wb_rf__T_120_data = 32'h0;
  assign wb_rf__T_120_addr = 5'h1d;
  assign wb_rf__T_120_mask = 1'h1;
  assign wb_rf__T_120_en = reset;
  assign wb_rf__T_124_data = 32'h0;
  assign wb_rf__T_124_addr = 5'h1e;
  assign wb_rf__T_124_mask = 1'h1;
  assign wb_rf__T_124_en = reset;
  assign wb_rf__T_128_data = 32'h0;
  assign wb_rf__T_128_addr = 5'h1f;
  assign wb_rf__T_128_mask = 1'h1;
  assign wb_rf__T_128_en = reset;
  assign wb_rf__T_182_data = io_wb_bits_data;
  assign wb_rf__T_182_addr = io_wb_bits_rd_idx;
  assign wb_rf__T_182_mask = 1'h1;
  assign wb_rf__T_182_en = _T_179 & _T_181;
  assign bp_rf__T_149_addr = io_rfio_rs_idx;
  assign bp_rf__T_149_data = bp_rf[bp_rf__T_149_addr]; // @[rf.scala 23:18]
  assign bp_rf__T_174_addr = io_rfio_rt_idx;
  assign bp_rf__T_174_data = bp_rf[bp_rf__T_174_addr]; // @[rf.scala 23:18]
  assign bp_rf__T_190_data = io_bp_bits_data;
  assign bp_rf__T_190_addr = io_bp_bits_rd_idx;
  assign bp_rf__T_190_mask = 1'h1;
  assign bp_rf__T_190_en = _T_134 & _T_188;
  assign rf_dirtys__T_129_addr = io_rfio_rs_idx;
  assign rf_dirtys__T_129_data = rf_dirtys[rf_dirtys__T_129_addr]; // @[rf.scala 24:22]
  assign rf_dirtys__T_141_addr = io_rfio_rs_idx;
  assign rf_dirtys__T_141_data = rf_dirtys[rf_dirtys__T_141_addr]; // @[rf.scala 24:22]
  assign rf_dirtys__T_154_addr = io_rfio_rt_idx;
  assign rf_dirtys__T_154_data = rf_dirtys[rf_dirtys__T_154_addr]; // @[rf.scala 24:22]
  assign rf_dirtys__T_166_addr = io_rfio_rt_idx;
  assign rf_dirtys__T_166_data = rf_dirtys[rf_dirtys__T_166_addr]; // @[rf.scala 24:22]
  assign rf_dirtys__T_2_data = 1'h0;
  assign rf_dirtys__T_2_addr = 5'h0;
  assign rf_dirtys__T_2_mask = 1'h1;
  assign rf_dirtys__T_2_en = reset;
  assign rf_dirtys__T_6_data = 1'h0;
  assign rf_dirtys__T_6_addr = 5'h1;
  assign rf_dirtys__T_6_mask = 1'h1;
  assign rf_dirtys__T_6_en = reset;
  assign rf_dirtys__T_10_data = 1'h0;
  assign rf_dirtys__T_10_addr = 5'h2;
  assign rf_dirtys__T_10_mask = 1'h1;
  assign rf_dirtys__T_10_en = reset;
  assign rf_dirtys__T_14_data = 1'h0;
  assign rf_dirtys__T_14_addr = 5'h3;
  assign rf_dirtys__T_14_mask = 1'h1;
  assign rf_dirtys__T_14_en = reset;
  assign rf_dirtys__T_18_data = 1'h0;
  assign rf_dirtys__T_18_addr = 5'h4;
  assign rf_dirtys__T_18_mask = 1'h1;
  assign rf_dirtys__T_18_en = reset;
  assign rf_dirtys__T_22_data = 1'h0;
  assign rf_dirtys__T_22_addr = 5'h5;
  assign rf_dirtys__T_22_mask = 1'h1;
  assign rf_dirtys__T_22_en = reset;
  assign rf_dirtys__T_26_data = 1'h0;
  assign rf_dirtys__T_26_addr = 5'h6;
  assign rf_dirtys__T_26_mask = 1'h1;
  assign rf_dirtys__T_26_en = reset;
  assign rf_dirtys__T_30_data = 1'h0;
  assign rf_dirtys__T_30_addr = 5'h7;
  assign rf_dirtys__T_30_mask = 1'h1;
  assign rf_dirtys__T_30_en = reset;
  assign rf_dirtys__T_34_data = 1'h0;
  assign rf_dirtys__T_34_addr = 5'h8;
  assign rf_dirtys__T_34_mask = 1'h1;
  assign rf_dirtys__T_34_en = reset;
  assign rf_dirtys__T_38_data = 1'h0;
  assign rf_dirtys__T_38_addr = 5'h9;
  assign rf_dirtys__T_38_mask = 1'h1;
  assign rf_dirtys__T_38_en = reset;
  assign rf_dirtys__T_42_data = 1'h0;
  assign rf_dirtys__T_42_addr = 5'ha;
  assign rf_dirtys__T_42_mask = 1'h1;
  assign rf_dirtys__T_42_en = reset;
  assign rf_dirtys__T_46_data = 1'h0;
  assign rf_dirtys__T_46_addr = 5'hb;
  assign rf_dirtys__T_46_mask = 1'h1;
  assign rf_dirtys__T_46_en = reset;
  assign rf_dirtys__T_50_data = 1'h0;
  assign rf_dirtys__T_50_addr = 5'hc;
  assign rf_dirtys__T_50_mask = 1'h1;
  assign rf_dirtys__T_50_en = reset;
  assign rf_dirtys__T_54_data = 1'h0;
  assign rf_dirtys__T_54_addr = 5'hd;
  assign rf_dirtys__T_54_mask = 1'h1;
  assign rf_dirtys__T_54_en = reset;
  assign rf_dirtys__T_58_data = 1'h0;
  assign rf_dirtys__T_58_addr = 5'he;
  assign rf_dirtys__T_58_mask = 1'h1;
  assign rf_dirtys__T_58_en = reset;
  assign rf_dirtys__T_62_data = 1'h0;
  assign rf_dirtys__T_62_addr = 5'hf;
  assign rf_dirtys__T_62_mask = 1'h1;
  assign rf_dirtys__T_62_en = reset;
  assign rf_dirtys__T_66_data = 1'h0;
  assign rf_dirtys__T_66_addr = 5'h10;
  assign rf_dirtys__T_66_mask = 1'h1;
  assign rf_dirtys__T_66_en = reset;
  assign rf_dirtys__T_70_data = 1'h0;
  assign rf_dirtys__T_70_addr = 5'h11;
  assign rf_dirtys__T_70_mask = 1'h1;
  assign rf_dirtys__T_70_en = reset;
  assign rf_dirtys__T_74_data = 1'h0;
  assign rf_dirtys__T_74_addr = 5'h12;
  assign rf_dirtys__T_74_mask = 1'h1;
  assign rf_dirtys__T_74_en = reset;
  assign rf_dirtys__T_78_data = 1'h0;
  assign rf_dirtys__T_78_addr = 5'h13;
  assign rf_dirtys__T_78_mask = 1'h1;
  assign rf_dirtys__T_78_en = reset;
  assign rf_dirtys__T_82_data = 1'h0;
  assign rf_dirtys__T_82_addr = 5'h14;
  assign rf_dirtys__T_82_mask = 1'h1;
  assign rf_dirtys__T_82_en = reset;
  assign rf_dirtys__T_86_data = 1'h0;
  assign rf_dirtys__T_86_addr = 5'h15;
  assign rf_dirtys__T_86_mask = 1'h1;
  assign rf_dirtys__T_86_en = reset;
  assign rf_dirtys__T_90_data = 1'h0;
  assign rf_dirtys__T_90_addr = 5'h16;
  assign rf_dirtys__T_90_mask = 1'h1;
  assign rf_dirtys__T_90_en = reset;
  assign rf_dirtys__T_94_data = 1'h0;
  assign rf_dirtys__T_94_addr = 5'h17;
  assign rf_dirtys__T_94_mask = 1'h1;
  assign rf_dirtys__T_94_en = reset;
  assign rf_dirtys__T_98_data = 1'h0;
  assign rf_dirtys__T_98_addr = 5'h18;
  assign rf_dirtys__T_98_mask = 1'h1;
  assign rf_dirtys__T_98_en = reset;
  assign rf_dirtys__T_102_data = 1'h0;
  assign rf_dirtys__T_102_addr = 5'h19;
  assign rf_dirtys__T_102_mask = 1'h1;
  assign rf_dirtys__T_102_en = reset;
  assign rf_dirtys__T_106_data = 1'h0;
  assign rf_dirtys__T_106_addr = 5'h1a;
  assign rf_dirtys__T_106_mask = 1'h1;
  assign rf_dirtys__T_106_en = reset;
  assign rf_dirtys__T_110_data = 1'h0;
  assign rf_dirtys__T_110_addr = 5'h1b;
  assign rf_dirtys__T_110_mask = 1'h1;
  assign rf_dirtys__T_110_en = reset;
  assign rf_dirtys__T_114_data = 1'h0;
  assign rf_dirtys__T_114_addr = 5'h1c;
  assign rf_dirtys__T_114_mask = 1'h1;
  assign rf_dirtys__T_114_en = reset;
  assign rf_dirtys__T_118_data = 1'h0;
  assign rf_dirtys__T_118_addr = 5'h1d;
  assign rf_dirtys__T_118_mask = 1'h1;
  assign rf_dirtys__T_118_en = reset;
  assign rf_dirtys__T_122_data = 1'h0;
  assign rf_dirtys__T_122_addr = 5'h1e;
  assign rf_dirtys__T_122_mask = 1'h1;
  assign rf_dirtys__T_122_en = reset;
  assign rf_dirtys__T_126_data = 1'h0;
  assign rf_dirtys__T_126_addr = 5'h1f;
  assign rf_dirtys__T_126_mask = 1'h1;
  assign rf_dirtys__T_126_en = reset;
  assign rf_dirtys__T_185_data = 1'h0;
  assign rf_dirtys__T_185_addr = io_wb_bits_rd_idx;
  assign rf_dirtys__T_185_mask = 1'h1;
  assign rf_dirtys__T_185_en = _T_179 & _T_184;
  assign rf_dirtys__T_192_data = 1'h1;
  assign rf_dirtys__T_192_addr = io_rfio_rd_idx;
  assign rf_dirtys__T_192_mask = 1'h1;
  assign rf_dirtys__T_192_en = io_rfio_wen;
  assign rf_dirtys__T_195_data = 1'h0;
  assign rf_dirtys__T_195_addr = 5'h0;
  assign rf_dirtys__T_195_mask = 1'h1;
  assign rf_dirtys__T_195_en = io_ex_flush_valid;
  assign rf_dirtys__T_197_data = 1'h0;
  assign rf_dirtys__T_197_addr = 5'h1;
  assign rf_dirtys__T_197_mask = 1'h1;
  assign rf_dirtys__T_197_en = io_ex_flush_valid;
  assign rf_dirtys__T_199_data = 1'h0;
  assign rf_dirtys__T_199_addr = 5'h2;
  assign rf_dirtys__T_199_mask = 1'h1;
  assign rf_dirtys__T_199_en = io_ex_flush_valid;
  assign rf_dirtys__T_201_data = 1'h0;
  assign rf_dirtys__T_201_addr = 5'h3;
  assign rf_dirtys__T_201_mask = 1'h1;
  assign rf_dirtys__T_201_en = io_ex_flush_valid;
  assign rf_dirtys__T_203_data = 1'h0;
  assign rf_dirtys__T_203_addr = 5'h4;
  assign rf_dirtys__T_203_mask = 1'h1;
  assign rf_dirtys__T_203_en = io_ex_flush_valid;
  assign rf_dirtys__T_205_data = 1'h0;
  assign rf_dirtys__T_205_addr = 5'h5;
  assign rf_dirtys__T_205_mask = 1'h1;
  assign rf_dirtys__T_205_en = io_ex_flush_valid;
  assign rf_dirtys__T_207_data = 1'h0;
  assign rf_dirtys__T_207_addr = 5'h6;
  assign rf_dirtys__T_207_mask = 1'h1;
  assign rf_dirtys__T_207_en = io_ex_flush_valid;
  assign rf_dirtys__T_209_data = 1'h0;
  assign rf_dirtys__T_209_addr = 5'h7;
  assign rf_dirtys__T_209_mask = 1'h1;
  assign rf_dirtys__T_209_en = io_ex_flush_valid;
  assign rf_dirtys__T_211_data = 1'h0;
  assign rf_dirtys__T_211_addr = 5'h8;
  assign rf_dirtys__T_211_mask = 1'h1;
  assign rf_dirtys__T_211_en = io_ex_flush_valid;
  assign rf_dirtys__T_213_data = 1'h0;
  assign rf_dirtys__T_213_addr = 5'h9;
  assign rf_dirtys__T_213_mask = 1'h1;
  assign rf_dirtys__T_213_en = io_ex_flush_valid;
  assign rf_dirtys__T_215_data = 1'h0;
  assign rf_dirtys__T_215_addr = 5'ha;
  assign rf_dirtys__T_215_mask = 1'h1;
  assign rf_dirtys__T_215_en = io_ex_flush_valid;
  assign rf_dirtys__T_217_data = 1'h0;
  assign rf_dirtys__T_217_addr = 5'hb;
  assign rf_dirtys__T_217_mask = 1'h1;
  assign rf_dirtys__T_217_en = io_ex_flush_valid;
  assign rf_dirtys__T_219_data = 1'h0;
  assign rf_dirtys__T_219_addr = 5'hc;
  assign rf_dirtys__T_219_mask = 1'h1;
  assign rf_dirtys__T_219_en = io_ex_flush_valid;
  assign rf_dirtys__T_221_data = 1'h0;
  assign rf_dirtys__T_221_addr = 5'hd;
  assign rf_dirtys__T_221_mask = 1'h1;
  assign rf_dirtys__T_221_en = io_ex_flush_valid;
  assign rf_dirtys__T_223_data = 1'h0;
  assign rf_dirtys__T_223_addr = 5'he;
  assign rf_dirtys__T_223_mask = 1'h1;
  assign rf_dirtys__T_223_en = io_ex_flush_valid;
  assign rf_dirtys__T_225_data = 1'h0;
  assign rf_dirtys__T_225_addr = 5'hf;
  assign rf_dirtys__T_225_mask = 1'h1;
  assign rf_dirtys__T_225_en = io_ex_flush_valid;
  assign rf_dirtys__T_227_data = 1'h0;
  assign rf_dirtys__T_227_addr = 5'h10;
  assign rf_dirtys__T_227_mask = 1'h1;
  assign rf_dirtys__T_227_en = io_ex_flush_valid;
  assign rf_dirtys__T_229_data = 1'h0;
  assign rf_dirtys__T_229_addr = 5'h11;
  assign rf_dirtys__T_229_mask = 1'h1;
  assign rf_dirtys__T_229_en = io_ex_flush_valid;
  assign rf_dirtys__T_231_data = 1'h0;
  assign rf_dirtys__T_231_addr = 5'h12;
  assign rf_dirtys__T_231_mask = 1'h1;
  assign rf_dirtys__T_231_en = io_ex_flush_valid;
  assign rf_dirtys__T_233_data = 1'h0;
  assign rf_dirtys__T_233_addr = 5'h13;
  assign rf_dirtys__T_233_mask = 1'h1;
  assign rf_dirtys__T_233_en = io_ex_flush_valid;
  assign rf_dirtys__T_235_data = 1'h0;
  assign rf_dirtys__T_235_addr = 5'h14;
  assign rf_dirtys__T_235_mask = 1'h1;
  assign rf_dirtys__T_235_en = io_ex_flush_valid;
  assign rf_dirtys__T_237_data = 1'h0;
  assign rf_dirtys__T_237_addr = 5'h15;
  assign rf_dirtys__T_237_mask = 1'h1;
  assign rf_dirtys__T_237_en = io_ex_flush_valid;
  assign rf_dirtys__T_239_data = 1'h0;
  assign rf_dirtys__T_239_addr = 5'h16;
  assign rf_dirtys__T_239_mask = 1'h1;
  assign rf_dirtys__T_239_en = io_ex_flush_valid;
  assign rf_dirtys__T_241_data = 1'h0;
  assign rf_dirtys__T_241_addr = 5'h17;
  assign rf_dirtys__T_241_mask = 1'h1;
  assign rf_dirtys__T_241_en = io_ex_flush_valid;
  assign rf_dirtys__T_243_data = 1'h0;
  assign rf_dirtys__T_243_addr = 5'h18;
  assign rf_dirtys__T_243_mask = 1'h1;
  assign rf_dirtys__T_243_en = io_ex_flush_valid;
  assign rf_dirtys__T_245_data = 1'h0;
  assign rf_dirtys__T_245_addr = 5'h19;
  assign rf_dirtys__T_245_mask = 1'h1;
  assign rf_dirtys__T_245_en = io_ex_flush_valid;
  assign rf_dirtys__T_247_data = 1'h0;
  assign rf_dirtys__T_247_addr = 5'h1a;
  assign rf_dirtys__T_247_mask = 1'h1;
  assign rf_dirtys__T_247_en = io_ex_flush_valid;
  assign rf_dirtys__T_249_data = 1'h0;
  assign rf_dirtys__T_249_addr = 5'h1b;
  assign rf_dirtys__T_249_mask = 1'h1;
  assign rf_dirtys__T_249_en = io_ex_flush_valid;
  assign rf_dirtys__T_251_data = 1'h0;
  assign rf_dirtys__T_251_addr = 5'h1c;
  assign rf_dirtys__T_251_mask = 1'h1;
  assign rf_dirtys__T_251_en = io_ex_flush_valid;
  assign rf_dirtys__T_253_data = 1'h0;
  assign rf_dirtys__T_253_addr = 5'h1d;
  assign rf_dirtys__T_253_mask = 1'h1;
  assign rf_dirtys__T_253_en = io_ex_flush_valid;
  assign rf_dirtys__T_255_data = 1'h0;
  assign rf_dirtys__T_255_addr = 5'h1e;
  assign rf_dirtys__T_255_mask = 1'h1;
  assign rf_dirtys__T_255_en = io_ex_flush_valid;
  assign rf_dirtys__T_257_data = 1'h0;
  assign rf_dirtys__T_257_addr = 5'h1f;
  assign rf_dirtys__T_257_mask = 1'h1;
  assign rf_dirtys__T_257_en = io_ex_flush_valid;
  assign bp_readys__T_131_addr = io_rfio_rs_idx;
  assign bp_readys__T_131_data = bp_readys[bp_readys__T_131_addr]; // @[rf.scala 25:22]
  assign bp_readys__T_148_addr = io_rfio_rs_idx;
  assign bp_readys__T_148_data = bp_readys[bp_readys__T_148_addr]; // @[rf.scala 25:22]
  assign bp_readys__T_156_addr = io_rfio_rt_idx;
  assign bp_readys__T_156_data = bp_readys[bp_readys__T_156_addr]; // @[rf.scala 25:22]
  assign bp_readys__T_173_addr = io_rfio_rt_idx;
  assign bp_readys__T_173_data = bp_readys[bp_readys__T_173_addr]; // @[rf.scala 25:22]
  assign bp_readys__T_3_data = 1'h0;
  assign bp_readys__T_3_addr = 5'h0;
  assign bp_readys__T_3_mask = 1'h1;
  assign bp_readys__T_3_en = reset;
  assign bp_readys__T_7_data = 1'h0;
  assign bp_readys__T_7_addr = 5'h1;
  assign bp_readys__T_7_mask = 1'h1;
  assign bp_readys__T_7_en = reset;
  assign bp_readys__T_11_data = 1'h0;
  assign bp_readys__T_11_addr = 5'h2;
  assign bp_readys__T_11_mask = 1'h1;
  assign bp_readys__T_11_en = reset;
  assign bp_readys__T_15_data = 1'h0;
  assign bp_readys__T_15_addr = 5'h3;
  assign bp_readys__T_15_mask = 1'h1;
  assign bp_readys__T_15_en = reset;
  assign bp_readys__T_19_data = 1'h0;
  assign bp_readys__T_19_addr = 5'h4;
  assign bp_readys__T_19_mask = 1'h1;
  assign bp_readys__T_19_en = reset;
  assign bp_readys__T_23_data = 1'h0;
  assign bp_readys__T_23_addr = 5'h5;
  assign bp_readys__T_23_mask = 1'h1;
  assign bp_readys__T_23_en = reset;
  assign bp_readys__T_27_data = 1'h0;
  assign bp_readys__T_27_addr = 5'h6;
  assign bp_readys__T_27_mask = 1'h1;
  assign bp_readys__T_27_en = reset;
  assign bp_readys__T_31_data = 1'h0;
  assign bp_readys__T_31_addr = 5'h7;
  assign bp_readys__T_31_mask = 1'h1;
  assign bp_readys__T_31_en = reset;
  assign bp_readys__T_35_data = 1'h0;
  assign bp_readys__T_35_addr = 5'h8;
  assign bp_readys__T_35_mask = 1'h1;
  assign bp_readys__T_35_en = reset;
  assign bp_readys__T_39_data = 1'h0;
  assign bp_readys__T_39_addr = 5'h9;
  assign bp_readys__T_39_mask = 1'h1;
  assign bp_readys__T_39_en = reset;
  assign bp_readys__T_43_data = 1'h0;
  assign bp_readys__T_43_addr = 5'ha;
  assign bp_readys__T_43_mask = 1'h1;
  assign bp_readys__T_43_en = reset;
  assign bp_readys__T_47_data = 1'h0;
  assign bp_readys__T_47_addr = 5'hb;
  assign bp_readys__T_47_mask = 1'h1;
  assign bp_readys__T_47_en = reset;
  assign bp_readys__T_51_data = 1'h0;
  assign bp_readys__T_51_addr = 5'hc;
  assign bp_readys__T_51_mask = 1'h1;
  assign bp_readys__T_51_en = reset;
  assign bp_readys__T_55_data = 1'h0;
  assign bp_readys__T_55_addr = 5'hd;
  assign bp_readys__T_55_mask = 1'h1;
  assign bp_readys__T_55_en = reset;
  assign bp_readys__T_59_data = 1'h0;
  assign bp_readys__T_59_addr = 5'he;
  assign bp_readys__T_59_mask = 1'h1;
  assign bp_readys__T_59_en = reset;
  assign bp_readys__T_63_data = 1'h0;
  assign bp_readys__T_63_addr = 5'hf;
  assign bp_readys__T_63_mask = 1'h1;
  assign bp_readys__T_63_en = reset;
  assign bp_readys__T_67_data = 1'h0;
  assign bp_readys__T_67_addr = 5'h10;
  assign bp_readys__T_67_mask = 1'h1;
  assign bp_readys__T_67_en = reset;
  assign bp_readys__T_71_data = 1'h0;
  assign bp_readys__T_71_addr = 5'h11;
  assign bp_readys__T_71_mask = 1'h1;
  assign bp_readys__T_71_en = reset;
  assign bp_readys__T_75_data = 1'h0;
  assign bp_readys__T_75_addr = 5'h12;
  assign bp_readys__T_75_mask = 1'h1;
  assign bp_readys__T_75_en = reset;
  assign bp_readys__T_79_data = 1'h0;
  assign bp_readys__T_79_addr = 5'h13;
  assign bp_readys__T_79_mask = 1'h1;
  assign bp_readys__T_79_en = reset;
  assign bp_readys__T_83_data = 1'h0;
  assign bp_readys__T_83_addr = 5'h14;
  assign bp_readys__T_83_mask = 1'h1;
  assign bp_readys__T_83_en = reset;
  assign bp_readys__T_87_data = 1'h0;
  assign bp_readys__T_87_addr = 5'h15;
  assign bp_readys__T_87_mask = 1'h1;
  assign bp_readys__T_87_en = reset;
  assign bp_readys__T_91_data = 1'h0;
  assign bp_readys__T_91_addr = 5'h16;
  assign bp_readys__T_91_mask = 1'h1;
  assign bp_readys__T_91_en = reset;
  assign bp_readys__T_95_data = 1'h0;
  assign bp_readys__T_95_addr = 5'h17;
  assign bp_readys__T_95_mask = 1'h1;
  assign bp_readys__T_95_en = reset;
  assign bp_readys__T_99_data = 1'h0;
  assign bp_readys__T_99_addr = 5'h18;
  assign bp_readys__T_99_mask = 1'h1;
  assign bp_readys__T_99_en = reset;
  assign bp_readys__T_103_data = 1'h0;
  assign bp_readys__T_103_addr = 5'h19;
  assign bp_readys__T_103_mask = 1'h1;
  assign bp_readys__T_103_en = reset;
  assign bp_readys__T_107_data = 1'h0;
  assign bp_readys__T_107_addr = 5'h1a;
  assign bp_readys__T_107_mask = 1'h1;
  assign bp_readys__T_107_en = reset;
  assign bp_readys__T_111_data = 1'h0;
  assign bp_readys__T_111_addr = 5'h1b;
  assign bp_readys__T_111_mask = 1'h1;
  assign bp_readys__T_111_en = reset;
  assign bp_readys__T_115_data = 1'h0;
  assign bp_readys__T_115_addr = 5'h1c;
  assign bp_readys__T_115_mask = 1'h1;
  assign bp_readys__T_115_en = reset;
  assign bp_readys__T_119_data = 1'h0;
  assign bp_readys__T_119_addr = 5'h1d;
  assign bp_readys__T_119_mask = 1'h1;
  assign bp_readys__T_119_en = reset;
  assign bp_readys__T_123_data = 1'h0;
  assign bp_readys__T_123_addr = 5'h1e;
  assign bp_readys__T_123_mask = 1'h1;
  assign bp_readys__T_123_en = reset;
  assign bp_readys__T_127_data = 1'h0;
  assign bp_readys__T_127_addr = 5'h1f;
  assign bp_readys__T_127_mask = 1'h1;
  assign bp_readys__T_127_en = reset;
  assign bp_readys__T_191_data = 1'h1;
  assign bp_readys__T_191_addr = io_bp_bits_rd_idx;
  assign bp_readys__T_191_mask = 1'h1;
  assign bp_readys__T_191_en = _T_134 & _T_188;
  assign bp_readys__T_193_data = 1'h0;
  assign bp_readys__T_193_addr = io_rfio_rd_idx;
  assign bp_readys__T_193_mask = 1'h1;
  assign bp_readys__T_193_en = io_rfio_wen;
  assign bp_readys__T_196_data = 1'h1;
  assign bp_readys__T_196_addr = 5'h0;
  assign bp_readys__T_196_mask = 1'h1;
  assign bp_readys__T_196_en = io_ex_flush_valid;
  assign bp_readys__T_198_data = 1'h1;
  assign bp_readys__T_198_addr = 5'h1;
  assign bp_readys__T_198_mask = 1'h1;
  assign bp_readys__T_198_en = io_ex_flush_valid;
  assign bp_readys__T_200_data = 1'h1;
  assign bp_readys__T_200_addr = 5'h2;
  assign bp_readys__T_200_mask = 1'h1;
  assign bp_readys__T_200_en = io_ex_flush_valid;
  assign bp_readys__T_202_data = 1'h1;
  assign bp_readys__T_202_addr = 5'h3;
  assign bp_readys__T_202_mask = 1'h1;
  assign bp_readys__T_202_en = io_ex_flush_valid;
  assign bp_readys__T_204_data = 1'h1;
  assign bp_readys__T_204_addr = 5'h4;
  assign bp_readys__T_204_mask = 1'h1;
  assign bp_readys__T_204_en = io_ex_flush_valid;
  assign bp_readys__T_206_data = 1'h1;
  assign bp_readys__T_206_addr = 5'h5;
  assign bp_readys__T_206_mask = 1'h1;
  assign bp_readys__T_206_en = io_ex_flush_valid;
  assign bp_readys__T_208_data = 1'h1;
  assign bp_readys__T_208_addr = 5'h6;
  assign bp_readys__T_208_mask = 1'h1;
  assign bp_readys__T_208_en = io_ex_flush_valid;
  assign bp_readys__T_210_data = 1'h1;
  assign bp_readys__T_210_addr = 5'h7;
  assign bp_readys__T_210_mask = 1'h1;
  assign bp_readys__T_210_en = io_ex_flush_valid;
  assign bp_readys__T_212_data = 1'h1;
  assign bp_readys__T_212_addr = 5'h8;
  assign bp_readys__T_212_mask = 1'h1;
  assign bp_readys__T_212_en = io_ex_flush_valid;
  assign bp_readys__T_214_data = 1'h1;
  assign bp_readys__T_214_addr = 5'h9;
  assign bp_readys__T_214_mask = 1'h1;
  assign bp_readys__T_214_en = io_ex_flush_valid;
  assign bp_readys__T_216_data = 1'h1;
  assign bp_readys__T_216_addr = 5'ha;
  assign bp_readys__T_216_mask = 1'h1;
  assign bp_readys__T_216_en = io_ex_flush_valid;
  assign bp_readys__T_218_data = 1'h1;
  assign bp_readys__T_218_addr = 5'hb;
  assign bp_readys__T_218_mask = 1'h1;
  assign bp_readys__T_218_en = io_ex_flush_valid;
  assign bp_readys__T_220_data = 1'h1;
  assign bp_readys__T_220_addr = 5'hc;
  assign bp_readys__T_220_mask = 1'h1;
  assign bp_readys__T_220_en = io_ex_flush_valid;
  assign bp_readys__T_222_data = 1'h1;
  assign bp_readys__T_222_addr = 5'hd;
  assign bp_readys__T_222_mask = 1'h1;
  assign bp_readys__T_222_en = io_ex_flush_valid;
  assign bp_readys__T_224_data = 1'h1;
  assign bp_readys__T_224_addr = 5'he;
  assign bp_readys__T_224_mask = 1'h1;
  assign bp_readys__T_224_en = io_ex_flush_valid;
  assign bp_readys__T_226_data = 1'h1;
  assign bp_readys__T_226_addr = 5'hf;
  assign bp_readys__T_226_mask = 1'h1;
  assign bp_readys__T_226_en = io_ex_flush_valid;
  assign bp_readys__T_228_data = 1'h1;
  assign bp_readys__T_228_addr = 5'h10;
  assign bp_readys__T_228_mask = 1'h1;
  assign bp_readys__T_228_en = io_ex_flush_valid;
  assign bp_readys__T_230_data = 1'h1;
  assign bp_readys__T_230_addr = 5'h11;
  assign bp_readys__T_230_mask = 1'h1;
  assign bp_readys__T_230_en = io_ex_flush_valid;
  assign bp_readys__T_232_data = 1'h1;
  assign bp_readys__T_232_addr = 5'h12;
  assign bp_readys__T_232_mask = 1'h1;
  assign bp_readys__T_232_en = io_ex_flush_valid;
  assign bp_readys__T_234_data = 1'h1;
  assign bp_readys__T_234_addr = 5'h13;
  assign bp_readys__T_234_mask = 1'h1;
  assign bp_readys__T_234_en = io_ex_flush_valid;
  assign bp_readys__T_236_data = 1'h1;
  assign bp_readys__T_236_addr = 5'h14;
  assign bp_readys__T_236_mask = 1'h1;
  assign bp_readys__T_236_en = io_ex_flush_valid;
  assign bp_readys__T_238_data = 1'h1;
  assign bp_readys__T_238_addr = 5'h15;
  assign bp_readys__T_238_mask = 1'h1;
  assign bp_readys__T_238_en = io_ex_flush_valid;
  assign bp_readys__T_240_data = 1'h1;
  assign bp_readys__T_240_addr = 5'h16;
  assign bp_readys__T_240_mask = 1'h1;
  assign bp_readys__T_240_en = io_ex_flush_valid;
  assign bp_readys__T_242_data = 1'h1;
  assign bp_readys__T_242_addr = 5'h17;
  assign bp_readys__T_242_mask = 1'h1;
  assign bp_readys__T_242_en = io_ex_flush_valid;
  assign bp_readys__T_244_data = 1'h1;
  assign bp_readys__T_244_addr = 5'h18;
  assign bp_readys__T_244_mask = 1'h1;
  assign bp_readys__T_244_en = io_ex_flush_valid;
  assign bp_readys__T_246_data = 1'h1;
  assign bp_readys__T_246_addr = 5'h19;
  assign bp_readys__T_246_mask = 1'h1;
  assign bp_readys__T_246_en = io_ex_flush_valid;
  assign bp_readys__T_248_data = 1'h1;
  assign bp_readys__T_248_addr = 5'h1a;
  assign bp_readys__T_248_mask = 1'h1;
  assign bp_readys__T_248_en = io_ex_flush_valid;
  assign bp_readys__T_250_data = 1'h1;
  assign bp_readys__T_250_addr = 5'h1b;
  assign bp_readys__T_250_mask = 1'h1;
  assign bp_readys__T_250_en = io_ex_flush_valid;
  assign bp_readys__T_252_data = 1'h1;
  assign bp_readys__T_252_addr = 5'h1c;
  assign bp_readys__T_252_mask = 1'h1;
  assign bp_readys__T_252_en = io_ex_flush_valid;
  assign bp_readys__T_254_data = 1'h1;
  assign bp_readys__T_254_addr = 5'h1d;
  assign bp_readys__T_254_mask = 1'h1;
  assign bp_readys__T_254_en = io_ex_flush_valid;
  assign bp_readys__T_256_data = 1'h1;
  assign bp_readys__T_256_addr = 5'h1e;
  assign bp_readys__T_256_mask = 1'h1;
  assign bp_readys__T_256_en = io_ex_flush_valid;
  assign bp_readys__T_258_data = 1'h1;
  assign bp_readys__T_258_addr = 5'h1f;
  assign bp_readys__T_258_mask = 1'h1;
  assign bp_readys__T_258_en = io_ex_flush_valid;
  assign io_rfio_rs_data_valid = _T_137 | _T_138; // @[rf.scala 44:25]
  assign io_rfio_rs_data_bits = _T_138 ? 32'h0 : _T_152; // @[rf.scala 45:24]
  assign io_rfio_rt_data_valid = _T_162 | _T_163; // @[rf.scala 47:25]
  assign io_rfio_rt_data_bits = _T_163 ? 32'h0 : _T_177; // @[rf.scala 48:24]
  assign io_commit_valid = io_wb_valid; // @[rf.scala 79:19]
  assign io_commit_pc = io_wb_bits_pc; // @[rf.scala 80:16]
  assign io_commit_instr = {_T_262,_T_260}; // @[rf.scala 81:19]
  assign io_commit_ip7 = io_wb_bits_ip7; // @[rf.scala 82:17]
  assign io_commit_gpr_0 = _T_267 ? io_wb_bits_data : wb_rf__T_268_data; // @[rf.scala 87:22]
  assign io_commit_gpr_1 = _T_272 ? io_wb_bits_data : wb_rf__T_273_data; // @[rf.scala 87:22]
  assign io_commit_gpr_2 = _T_277 ? io_wb_bits_data : wb_rf__T_278_data; // @[rf.scala 87:22]
  assign io_commit_gpr_3 = _T_282 ? io_wb_bits_data : wb_rf__T_283_data; // @[rf.scala 87:22]
  assign io_commit_gpr_4 = _T_287 ? io_wb_bits_data : wb_rf__T_288_data; // @[rf.scala 87:22]
  assign io_commit_gpr_5 = _T_292 ? io_wb_bits_data : wb_rf__T_293_data; // @[rf.scala 87:22]
  assign io_commit_gpr_6 = _T_297 ? io_wb_bits_data : wb_rf__T_298_data; // @[rf.scala 87:22]
  assign io_commit_gpr_7 = _T_302 ? io_wb_bits_data : wb_rf__T_303_data; // @[rf.scala 87:22]
  assign io_commit_gpr_8 = _T_307 ? io_wb_bits_data : wb_rf__T_308_data; // @[rf.scala 87:22]
  assign io_commit_gpr_9 = _T_312 ? io_wb_bits_data : wb_rf__T_313_data; // @[rf.scala 87:22]
  assign io_commit_gpr_10 = _T_317 ? io_wb_bits_data : wb_rf__T_318_data; // @[rf.scala 87:22]
  assign io_commit_gpr_11 = _T_322 ? io_wb_bits_data : wb_rf__T_323_data; // @[rf.scala 87:22]
  assign io_commit_gpr_12 = _T_327 ? io_wb_bits_data : wb_rf__T_328_data; // @[rf.scala 87:22]
  assign io_commit_gpr_13 = _T_332 ? io_wb_bits_data : wb_rf__T_333_data; // @[rf.scala 87:22]
  assign io_commit_gpr_14 = _T_337 ? io_wb_bits_data : wb_rf__T_338_data; // @[rf.scala 87:22]
  assign io_commit_gpr_15 = _T_342 ? io_wb_bits_data : wb_rf__T_343_data; // @[rf.scala 87:22]
  assign io_commit_gpr_16 = _T_347 ? io_wb_bits_data : wb_rf__T_348_data; // @[rf.scala 87:22]
  assign io_commit_gpr_17 = _T_352 ? io_wb_bits_data : wb_rf__T_353_data; // @[rf.scala 87:22]
  assign io_commit_gpr_18 = _T_357 ? io_wb_bits_data : wb_rf__T_358_data; // @[rf.scala 87:22]
  assign io_commit_gpr_19 = _T_362 ? io_wb_bits_data : wb_rf__T_363_data; // @[rf.scala 87:22]
  assign io_commit_gpr_20 = _T_367 ? io_wb_bits_data : wb_rf__T_368_data; // @[rf.scala 87:22]
  assign io_commit_gpr_21 = _T_372 ? io_wb_bits_data : wb_rf__T_373_data; // @[rf.scala 87:22]
  assign io_commit_gpr_22 = _T_377 ? io_wb_bits_data : wb_rf__T_378_data; // @[rf.scala 87:22]
  assign io_commit_gpr_23 = _T_382 ? io_wb_bits_data : wb_rf__T_383_data; // @[rf.scala 87:22]
  assign io_commit_gpr_24 = _T_387 ? io_wb_bits_data : wb_rf__T_388_data; // @[rf.scala 87:22]
  assign io_commit_gpr_25 = _T_392 ? io_wb_bits_data : wb_rf__T_393_data; // @[rf.scala 87:22]
  assign io_commit_gpr_26 = _T_397 ? io_wb_bits_data : wb_rf__T_398_data; // @[rf.scala 87:22]
  assign io_commit_gpr_27 = _T_402 ? io_wb_bits_data : wb_rf__T_403_data; // @[rf.scala 87:22]
  assign io_commit_gpr_28 = _T_407 ? io_wb_bits_data : wb_rf__T_408_data; // @[rf.scala 87:22]
  assign io_commit_gpr_29 = _T_412 ? io_wb_bits_data : wb_rf__T_413_data; // @[rf.scala 87:22]
  assign io_commit_gpr_30 = _T_417 ? io_wb_bits_data : wb_rf__T_418_data; // @[rf.scala 87:22]
  assign io_commit_gpr_31 = _T_422 ? io_wb_bits_data : wb_rf__T_423_data; // @[rf.scala 87:22]
  assign io_commit_rd_idx = io_wb_bits_rd_idx; // @[rf.scala 85:20]
  assign io_commit_wdata = io_wb_bits_data; // @[rf.scala 84:19]
  assign io_commit_wen = io_wb_bits_v & io_wb_bits_wen; // @[rf.scala 83:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    wbids[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    wb_rf[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    bp_rf[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rf_dirtys[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    bp_readys[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(wbids__T_1_en & wbids__T_1_mask) begin
      wbids[wbids__T_1_addr] <= wbids__T_1_data; // @[rf.scala 21:18]
    end
    if(wbids__T_5_en & wbids__T_5_mask) begin
      wbids[wbids__T_5_addr] <= wbids__T_5_data; // @[rf.scala 21:18]
    end
    if(wbids__T_9_en & wbids__T_9_mask) begin
      wbids[wbids__T_9_addr] <= wbids__T_9_data; // @[rf.scala 21:18]
    end
    if(wbids__T_13_en & wbids__T_13_mask) begin
      wbids[wbids__T_13_addr] <= wbids__T_13_data; // @[rf.scala 21:18]
    end
    if(wbids__T_17_en & wbids__T_17_mask) begin
      wbids[wbids__T_17_addr] <= wbids__T_17_data; // @[rf.scala 21:18]
    end
    if(wbids__T_21_en & wbids__T_21_mask) begin
      wbids[wbids__T_21_addr] <= wbids__T_21_data; // @[rf.scala 21:18]
    end
    if(wbids__T_25_en & wbids__T_25_mask) begin
      wbids[wbids__T_25_addr] <= wbids__T_25_data; // @[rf.scala 21:18]
    end
    if(wbids__T_29_en & wbids__T_29_mask) begin
      wbids[wbids__T_29_addr] <= wbids__T_29_data; // @[rf.scala 21:18]
    end
    if(wbids__T_33_en & wbids__T_33_mask) begin
      wbids[wbids__T_33_addr] <= wbids__T_33_data; // @[rf.scala 21:18]
    end
    if(wbids__T_37_en & wbids__T_37_mask) begin
      wbids[wbids__T_37_addr] <= wbids__T_37_data; // @[rf.scala 21:18]
    end
    if(wbids__T_41_en & wbids__T_41_mask) begin
      wbids[wbids__T_41_addr] <= wbids__T_41_data; // @[rf.scala 21:18]
    end
    if(wbids__T_45_en & wbids__T_45_mask) begin
      wbids[wbids__T_45_addr] <= wbids__T_45_data; // @[rf.scala 21:18]
    end
    if(wbids__T_49_en & wbids__T_49_mask) begin
      wbids[wbids__T_49_addr] <= wbids__T_49_data; // @[rf.scala 21:18]
    end
    if(wbids__T_53_en & wbids__T_53_mask) begin
      wbids[wbids__T_53_addr] <= wbids__T_53_data; // @[rf.scala 21:18]
    end
    if(wbids__T_57_en & wbids__T_57_mask) begin
      wbids[wbids__T_57_addr] <= wbids__T_57_data; // @[rf.scala 21:18]
    end
    if(wbids__T_61_en & wbids__T_61_mask) begin
      wbids[wbids__T_61_addr] <= wbids__T_61_data; // @[rf.scala 21:18]
    end
    if(wbids__T_65_en & wbids__T_65_mask) begin
      wbids[wbids__T_65_addr] <= wbids__T_65_data; // @[rf.scala 21:18]
    end
    if(wbids__T_69_en & wbids__T_69_mask) begin
      wbids[wbids__T_69_addr] <= wbids__T_69_data; // @[rf.scala 21:18]
    end
    if(wbids__T_73_en & wbids__T_73_mask) begin
      wbids[wbids__T_73_addr] <= wbids__T_73_data; // @[rf.scala 21:18]
    end
    if(wbids__T_77_en & wbids__T_77_mask) begin
      wbids[wbids__T_77_addr] <= wbids__T_77_data; // @[rf.scala 21:18]
    end
    if(wbids__T_81_en & wbids__T_81_mask) begin
      wbids[wbids__T_81_addr] <= wbids__T_81_data; // @[rf.scala 21:18]
    end
    if(wbids__T_85_en & wbids__T_85_mask) begin
      wbids[wbids__T_85_addr] <= wbids__T_85_data; // @[rf.scala 21:18]
    end
    if(wbids__T_89_en & wbids__T_89_mask) begin
      wbids[wbids__T_89_addr] <= wbids__T_89_data; // @[rf.scala 21:18]
    end
    if(wbids__T_93_en & wbids__T_93_mask) begin
      wbids[wbids__T_93_addr] <= wbids__T_93_data; // @[rf.scala 21:18]
    end
    if(wbids__T_97_en & wbids__T_97_mask) begin
      wbids[wbids__T_97_addr] <= wbids__T_97_data; // @[rf.scala 21:18]
    end
    if(wbids__T_101_en & wbids__T_101_mask) begin
      wbids[wbids__T_101_addr] <= wbids__T_101_data; // @[rf.scala 21:18]
    end
    if(wbids__T_105_en & wbids__T_105_mask) begin
      wbids[wbids__T_105_addr] <= wbids__T_105_data; // @[rf.scala 21:18]
    end
    if(wbids__T_109_en & wbids__T_109_mask) begin
      wbids[wbids__T_109_addr] <= wbids__T_109_data; // @[rf.scala 21:18]
    end
    if(wbids__T_113_en & wbids__T_113_mask) begin
      wbids[wbids__T_113_addr] <= wbids__T_113_data; // @[rf.scala 21:18]
    end
    if(wbids__T_117_en & wbids__T_117_mask) begin
      wbids[wbids__T_117_addr] <= wbids__T_117_data; // @[rf.scala 21:18]
    end
    if(wbids__T_121_en & wbids__T_121_mask) begin
      wbids[wbids__T_121_addr] <= wbids__T_121_data; // @[rf.scala 21:18]
    end
    if(wbids__T_125_en & wbids__T_125_mask) begin
      wbids[wbids__T_125_addr] <= wbids__T_125_data; // @[rf.scala 21:18]
    end
    if(wbids__T_194_en & wbids__T_194_mask) begin
      wbids[wbids__T_194_addr] <= wbids__T_194_data; // @[rf.scala 21:18]
    end
    if(wb_rf__T_4_en & wb_rf__T_4_mask) begin
      wb_rf[wb_rf__T_4_addr] <= wb_rf__T_4_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_8_en & wb_rf__T_8_mask) begin
      wb_rf[wb_rf__T_8_addr] <= wb_rf__T_8_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_12_en & wb_rf__T_12_mask) begin
      wb_rf[wb_rf__T_12_addr] <= wb_rf__T_12_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_16_en & wb_rf__T_16_mask) begin
      wb_rf[wb_rf__T_16_addr] <= wb_rf__T_16_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_20_en & wb_rf__T_20_mask) begin
      wb_rf[wb_rf__T_20_addr] <= wb_rf__T_20_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_24_en & wb_rf__T_24_mask) begin
      wb_rf[wb_rf__T_24_addr] <= wb_rf__T_24_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_28_en & wb_rf__T_28_mask) begin
      wb_rf[wb_rf__T_28_addr] <= wb_rf__T_28_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_32_en & wb_rf__T_32_mask) begin
      wb_rf[wb_rf__T_32_addr] <= wb_rf__T_32_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_36_en & wb_rf__T_36_mask) begin
      wb_rf[wb_rf__T_36_addr] <= wb_rf__T_36_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_40_en & wb_rf__T_40_mask) begin
      wb_rf[wb_rf__T_40_addr] <= wb_rf__T_40_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_44_en & wb_rf__T_44_mask) begin
      wb_rf[wb_rf__T_44_addr] <= wb_rf__T_44_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_48_en & wb_rf__T_48_mask) begin
      wb_rf[wb_rf__T_48_addr] <= wb_rf__T_48_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_52_en & wb_rf__T_52_mask) begin
      wb_rf[wb_rf__T_52_addr] <= wb_rf__T_52_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_56_en & wb_rf__T_56_mask) begin
      wb_rf[wb_rf__T_56_addr] <= wb_rf__T_56_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_60_en & wb_rf__T_60_mask) begin
      wb_rf[wb_rf__T_60_addr] <= wb_rf__T_60_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_64_en & wb_rf__T_64_mask) begin
      wb_rf[wb_rf__T_64_addr] <= wb_rf__T_64_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_68_en & wb_rf__T_68_mask) begin
      wb_rf[wb_rf__T_68_addr] <= wb_rf__T_68_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_72_en & wb_rf__T_72_mask) begin
      wb_rf[wb_rf__T_72_addr] <= wb_rf__T_72_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_76_en & wb_rf__T_76_mask) begin
      wb_rf[wb_rf__T_76_addr] <= wb_rf__T_76_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_80_en & wb_rf__T_80_mask) begin
      wb_rf[wb_rf__T_80_addr] <= wb_rf__T_80_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_84_en & wb_rf__T_84_mask) begin
      wb_rf[wb_rf__T_84_addr] <= wb_rf__T_84_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_88_en & wb_rf__T_88_mask) begin
      wb_rf[wb_rf__T_88_addr] <= wb_rf__T_88_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_92_en & wb_rf__T_92_mask) begin
      wb_rf[wb_rf__T_92_addr] <= wb_rf__T_92_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_96_en & wb_rf__T_96_mask) begin
      wb_rf[wb_rf__T_96_addr] <= wb_rf__T_96_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_100_en & wb_rf__T_100_mask) begin
      wb_rf[wb_rf__T_100_addr] <= wb_rf__T_100_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_104_en & wb_rf__T_104_mask) begin
      wb_rf[wb_rf__T_104_addr] <= wb_rf__T_104_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_108_en & wb_rf__T_108_mask) begin
      wb_rf[wb_rf__T_108_addr] <= wb_rf__T_108_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_112_en & wb_rf__T_112_mask) begin
      wb_rf[wb_rf__T_112_addr] <= wb_rf__T_112_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_116_en & wb_rf__T_116_mask) begin
      wb_rf[wb_rf__T_116_addr] <= wb_rf__T_116_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_120_en & wb_rf__T_120_mask) begin
      wb_rf[wb_rf__T_120_addr] <= wb_rf__T_120_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_124_en & wb_rf__T_124_mask) begin
      wb_rf[wb_rf__T_124_addr] <= wb_rf__T_124_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_128_en & wb_rf__T_128_mask) begin
      wb_rf[wb_rf__T_128_addr] <= wb_rf__T_128_data; // @[rf.scala 22:18]
    end
    if(wb_rf__T_182_en & wb_rf__T_182_mask) begin
      wb_rf[wb_rf__T_182_addr] <= wb_rf__T_182_data; // @[rf.scala 22:18]
    end
    if(bp_rf__T_190_en & bp_rf__T_190_mask) begin
      bp_rf[bp_rf__T_190_addr] <= bp_rf__T_190_data; // @[rf.scala 23:18]
    end
    if(rf_dirtys__T_2_en & rf_dirtys__T_2_mask) begin
      rf_dirtys[rf_dirtys__T_2_addr] <= rf_dirtys__T_2_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_6_en & rf_dirtys__T_6_mask) begin
      rf_dirtys[rf_dirtys__T_6_addr] <= rf_dirtys__T_6_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_10_en & rf_dirtys__T_10_mask) begin
      rf_dirtys[rf_dirtys__T_10_addr] <= rf_dirtys__T_10_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_14_en & rf_dirtys__T_14_mask) begin
      rf_dirtys[rf_dirtys__T_14_addr] <= rf_dirtys__T_14_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_18_en & rf_dirtys__T_18_mask) begin
      rf_dirtys[rf_dirtys__T_18_addr] <= rf_dirtys__T_18_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_22_en & rf_dirtys__T_22_mask) begin
      rf_dirtys[rf_dirtys__T_22_addr] <= rf_dirtys__T_22_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_26_en & rf_dirtys__T_26_mask) begin
      rf_dirtys[rf_dirtys__T_26_addr] <= rf_dirtys__T_26_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_30_en & rf_dirtys__T_30_mask) begin
      rf_dirtys[rf_dirtys__T_30_addr] <= rf_dirtys__T_30_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_34_en & rf_dirtys__T_34_mask) begin
      rf_dirtys[rf_dirtys__T_34_addr] <= rf_dirtys__T_34_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_38_en & rf_dirtys__T_38_mask) begin
      rf_dirtys[rf_dirtys__T_38_addr] <= rf_dirtys__T_38_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_42_en & rf_dirtys__T_42_mask) begin
      rf_dirtys[rf_dirtys__T_42_addr] <= rf_dirtys__T_42_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_46_en & rf_dirtys__T_46_mask) begin
      rf_dirtys[rf_dirtys__T_46_addr] <= rf_dirtys__T_46_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_50_en & rf_dirtys__T_50_mask) begin
      rf_dirtys[rf_dirtys__T_50_addr] <= rf_dirtys__T_50_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_54_en & rf_dirtys__T_54_mask) begin
      rf_dirtys[rf_dirtys__T_54_addr] <= rf_dirtys__T_54_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_58_en & rf_dirtys__T_58_mask) begin
      rf_dirtys[rf_dirtys__T_58_addr] <= rf_dirtys__T_58_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_62_en & rf_dirtys__T_62_mask) begin
      rf_dirtys[rf_dirtys__T_62_addr] <= rf_dirtys__T_62_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_66_en & rf_dirtys__T_66_mask) begin
      rf_dirtys[rf_dirtys__T_66_addr] <= rf_dirtys__T_66_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_70_en & rf_dirtys__T_70_mask) begin
      rf_dirtys[rf_dirtys__T_70_addr] <= rf_dirtys__T_70_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_74_en & rf_dirtys__T_74_mask) begin
      rf_dirtys[rf_dirtys__T_74_addr] <= rf_dirtys__T_74_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_78_en & rf_dirtys__T_78_mask) begin
      rf_dirtys[rf_dirtys__T_78_addr] <= rf_dirtys__T_78_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_82_en & rf_dirtys__T_82_mask) begin
      rf_dirtys[rf_dirtys__T_82_addr] <= rf_dirtys__T_82_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_86_en & rf_dirtys__T_86_mask) begin
      rf_dirtys[rf_dirtys__T_86_addr] <= rf_dirtys__T_86_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_90_en & rf_dirtys__T_90_mask) begin
      rf_dirtys[rf_dirtys__T_90_addr] <= rf_dirtys__T_90_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_94_en & rf_dirtys__T_94_mask) begin
      rf_dirtys[rf_dirtys__T_94_addr] <= rf_dirtys__T_94_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_98_en & rf_dirtys__T_98_mask) begin
      rf_dirtys[rf_dirtys__T_98_addr] <= rf_dirtys__T_98_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_102_en & rf_dirtys__T_102_mask) begin
      rf_dirtys[rf_dirtys__T_102_addr] <= rf_dirtys__T_102_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_106_en & rf_dirtys__T_106_mask) begin
      rf_dirtys[rf_dirtys__T_106_addr] <= rf_dirtys__T_106_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_110_en & rf_dirtys__T_110_mask) begin
      rf_dirtys[rf_dirtys__T_110_addr] <= rf_dirtys__T_110_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_114_en & rf_dirtys__T_114_mask) begin
      rf_dirtys[rf_dirtys__T_114_addr] <= rf_dirtys__T_114_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_118_en & rf_dirtys__T_118_mask) begin
      rf_dirtys[rf_dirtys__T_118_addr] <= rf_dirtys__T_118_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_122_en & rf_dirtys__T_122_mask) begin
      rf_dirtys[rf_dirtys__T_122_addr] <= rf_dirtys__T_122_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_126_en & rf_dirtys__T_126_mask) begin
      rf_dirtys[rf_dirtys__T_126_addr] <= rf_dirtys__T_126_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_185_en & rf_dirtys__T_185_mask) begin
      rf_dirtys[rf_dirtys__T_185_addr] <= rf_dirtys__T_185_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_192_en & rf_dirtys__T_192_mask) begin
      rf_dirtys[rf_dirtys__T_192_addr] <= rf_dirtys__T_192_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_195_en & rf_dirtys__T_195_mask) begin
      rf_dirtys[rf_dirtys__T_195_addr] <= rf_dirtys__T_195_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_197_en & rf_dirtys__T_197_mask) begin
      rf_dirtys[rf_dirtys__T_197_addr] <= rf_dirtys__T_197_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_199_en & rf_dirtys__T_199_mask) begin
      rf_dirtys[rf_dirtys__T_199_addr] <= rf_dirtys__T_199_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_201_en & rf_dirtys__T_201_mask) begin
      rf_dirtys[rf_dirtys__T_201_addr] <= rf_dirtys__T_201_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_203_en & rf_dirtys__T_203_mask) begin
      rf_dirtys[rf_dirtys__T_203_addr] <= rf_dirtys__T_203_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_205_en & rf_dirtys__T_205_mask) begin
      rf_dirtys[rf_dirtys__T_205_addr] <= rf_dirtys__T_205_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_207_en & rf_dirtys__T_207_mask) begin
      rf_dirtys[rf_dirtys__T_207_addr] <= rf_dirtys__T_207_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_209_en & rf_dirtys__T_209_mask) begin
      rf_dirtys[rf_dirtys__T_209_addr] <= rf_dirtys__T_209_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_211_en & rf_dirtys__T_211_mask) begin
      rf_dirtys[rf_dirtys__T_211_addr] <= rf_dirtys__T_211_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_213_en & rf_dirtys__T_213_mask) begin
      rf_dirtys[rf_dirtys__T_213_addr] <= rf_dirtys__T_213_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_215_en & rf_dirtys__T_215_mask) begin
      rf_dirtys[rf_dirtys__T_215_addr] <= rf_dirtys__T_215_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_217_en & rf_dirtys__T_217_mask) begin
      rf_dirtys[rf_dirtys__T_217_addr] <= rf_dirtys__T_217_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_219_en & rf_dirtys__T_219_mask) begin
      rf_dirtys[rf_dirtys__T_219_addr] <= rf_dirtys__T_219_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_221_en & rf_dirtys__T_221_mask) begin
      rf_dirtys[rf_dirtys__T_221_addr] <= rf_dirtys__T_221_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_223_en & rf_dirtys__T_223_mask) begin
      rf_dirtys[rf_dirtys__T_223_addr] <= rf_dirtys__T_223_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_225_en & rf_dirtys__T_225_mask) begin
      rf_dirtys[rf_dirtys__T_225_addr] <= rf_dirtys__T_225_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_227_en & rf_dirtys__T_227_mask) begin
      rf_dirtys[rf_dirtys__T_227_addr] <= rf_dirtys__T_227_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_229_en & rf_dirtys__T_229_mask) begin
      rf_dirtys[rf_dirtys__T_229_addr] <= rf_dirtys__T_229_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_231_en & rf_dirtys__T_231_mask) begin
      rf_dirtys[rf_dirtys__T_231_addr] <= rf_dirtys__T_231_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_233_en & rf_dirtys__T_233_mask) begin
      rf_dirtys[rf_dirtys__T_233_addr] <= rf_dirtys__T_233_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_235_en & rf_dirtys__T_235_mask) begin
      rf_dirtys[rf_dirtys__T_235_addr] <= rf_dirtys__T_235_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_237_en & rf_dirtys__T_237_mask) begin
      rf_dirtys[rf_dirtys__T_237_addr] <= rf_dirtys__T_237_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_239_en & rf_dirtys__T_239_mask) begin
      rf_dirtys[rf_dirtys__T_239_addr] <= rf_dirtys__T_239_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_241_en & rf_dirtys__T_241_mask) begin
      rf_dirtys[rf_dirtys__T_241_addr] <= rf_dirtys__T_241_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_243_en & rf_dirtys__T_243_mask) begin
      rf_dirtys[rf_dirtys__T_243_addr] <= rf_dirtys__T_243_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_245_en & rf_dirtys__T_245_mask) begin
      rf_dirtys[rf_dirtys__T_245_addr] <= rf_dirtys__T_245_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_247_en & rf_dirtys__T_247_mask) begin
      rf_dirtys[rf_dirtys__T_247_addr] <= rf_dirtys__T_247_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_249_en & rf_dirtys__T_249_mask) begin
      rf_dirtys[rf_dirtys__T_249_addr] <= rf_dirtys__T_249_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_251_en & rf_dirtys__T_251_mask) begin
      rf_dirtys[rf_dirtys__T_251_addr] <= rf_dirtys__T_251_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_253_en & rf_dirtys__T_253_mask) begin
      rf_dirtys[rf_dirtys__T_253_addr] <= rf_dirtys__T_253_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_255_en & rf_dirtys__T_255_mask) begin
      rf_dirtys[rf_dirtys__T_255_addr] <= rf_dirtys__T_255_data; // @[rf.scala 24:22]
    end
    if(rf_dirtys__T_257_en & rf_dirtys__T_257_mask) begin
      rf_dirtys[rf_dirtys__T_257_addr] <= rf_dirtys__T_257_data; // @[rf.scala 24:22]
    end
    if(bp_readys__T_3_en & bp_readys__T_3_mask) begin
      bp_readys[bp_readys__T_3_addr] <= bp_readys__T_3_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_7_en & bp_readys__T_7_mask) begin
      bp_readys[bp_readys__T_7_addr] <= bp_readys__T_7_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_11_en & bp_readys__T_11_mask) begin
      bp_readys[bp_readys__T_11_addr] <= bp_readys__T_11_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_15_en & bp_readys__T_15_mask) begin
      bp_readys[bp_readys__T_15_addr] <= bp_readys__T_15_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_19_en & bp_readys__T_19_mask) begin
      bp_readys[bp_readys__T_19_addr] <= bp_readys__T_19_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_23_en & bp_readys__T_23_mask) begin
      bp_readys[bp_readys__T_23_addr] <= bp_readys__T_23_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_27_en & bp_readys__T_27_mask) begin
      bp_readys[bp_readys__T_27_addr] <= bp_readys__T_27_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_31_en & bp_readys__T_31_mask) begin
      bp_readys[bp_readys__T_31_addr] <= bp_readys__T_31_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_35_en & bp_readys__T_35_mask) begin
      bp_readys[bp_readys__T_35_addr] <= bp_readys__T_35_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_39_en & bp_readys__T_39_mask) begin
      bp_readys[bp_readys__T_39_addr] <= bp_readys__T_39_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_43_en & bp_readys__T_43_mask) begin
      bp_readys[bp_readys__T_43_addr] <= bp_readys__T_43_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_47_en & bp_readys__T_47_mask) begin
      bp_readys[bp_readys__T_47_addr] <= bp_readys__T_47_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_51_en & bp_readys__T_51_mask) begin
      bp_readys[bp_readys__T_51_addr] <= bp_readys__T_51_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_55_en & bp_readys__T_55_mask) begin
      bp_readys[bp_readys__T_55_addr] <= bp_readys__T_55_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_59_en & bp_readys__T_59_mask) begin
      bp_readys[bp_readys__T_59_addr] <= bp_readys__T_59_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_63_en & bp_readys__T_63_mask) begin
      bp_readys[bp_readys__T_63_addr] <= bp_readys__T_63_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_67_en & bp_readys__T_67_mask) begin
      bp_readys[bp_readys__T_67_addr] <= bp_readys__T_67_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_71_en & bp_readys__T_71_mask) begin
      bp_readys[bp_readys__T_71_addr] <= bp_readys__T_71_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_75_en & bp_readys__T_75_mask) begin
      bp_readys[bp_readys__T_75_addr] <= bp_readys__T_75_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_79_en & bp_readys__T_79_mask) begin
      bp_readys[bp_readys__T_79_addr] <= bp_readys__T_79_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_83_en & bp_readys__T_83_mask) begin
      bp_readys[bp_readys__T_83_addr] <= bp_readys__T_83_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_87_en & bp_readys__T_87_mask) begin
      bp_readys[bp_readys__T_87_addr] <= bp_readys__T_87_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_91_en & bp_readys__T_91_mask) begin
      bp_readys[bp_readys__T_91_addr] <= bp_readys__T_91_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_95_en & bp_readys__T_95_mask) begin
      bp_readys[bp_readys__T_95_addr] <= bp_readys__T_95_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_99_en & bp_readys__T_99_mask) begin
      bp_readys[bp_readys__T_99_addr] <= bp_readys__T_99_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_103_en & bp_readys__T_103_mask) begin
      bp_readys[bp_readys__T_103_addr] <= bp_readys__T_103_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_107_en & bp_readys__T_107_mask) begin
      bp_readys[bp_readys__T_107_addr] <= bp_readys__T_107_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_111_en & bp_readys__T_111_mask) begin
      bp_readys[bp_readys__T_111_addr] <= bp_readys__T_111_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_115_en & bp_readys__T_115_mask) begin
      bp_readys[bp_readys__T_115_addr] <= bp_readys__T_115_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_119_en & bp_readys__T_119_mask) begin
      bp_readys[bp_readys__T_119_addr] <= bp_readys__T_119_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_123_en & bp_readys__T_123_mask) begin
      bp_readys[bp_readys__T_123_addr] <= bp_readys__T_123_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_127_en & bp_readys__T_127_mask) begin
      bp_readys[bp_readys__T_127_addr] <= bp_readys__T_127_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_191_en & bp_readys__T_191_mask) begin
      bp_readys[bp_readys__T_191_addr] <= bp_readys__T_191_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_193_en & bp_readys__T_193_mask) begin
      bp_readys[bp_readys__T_193_addr] <= bp_readys__T_193_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_196_en & bp_readys__T_196_mask) begin
      bp_readys[bp_readys__T_196_addr] <= bp_readys__T_196_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_198_en & bp_readys__T_198_mask) begin
      bp_readys[bp_readys__T_198_addr] <= bp_readys__T_198_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_200_en & bp_readys__T_200_mask) begin
      bp_readys[bp_readys__T_200_addr] <= bp_readys__T_200_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_202_en & bp_readys__T_202_mask) begin
      bp_readys[bp_readys__T_202_addr] <= bp_readys__T_202_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_204_en & bp_readys__T_204_mask) begin
      bp_readys[bp_readys__T_204_addr] <= bp_readys__T_204_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_206_en & bp_readys__T_206_mask) begin
      bp_readys[bp_readys__T_206_addr] <= bp_readys__T_206_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_208_en & bp_readys__T_208_mask) begin
      bp_readys[bp_readys__T_208_addr] <= bp_readys__T_208_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_210_en & bp_readys__T_210_mask) begin
      bp_readys[bp_readys__T_210_addr] <= bp_readys__T_210_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_212_en & bp_readys__T_212_mask) begin
      bp_readys[bp_readys__T_212_addr] <= bp_readys__T_212_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_214_en & bp_readys__T_214_mask) begin
      bp_readys[bp_readys__T_214_addr] <= bp_readys__T_214_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_216_en & bp_readys__T_216_mask) begin
      bp_readys[bp_readys__T_216_addr] <= bp_readys__T_216_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_218_en & bp_readys__T_218_mask) begin
      bp_readys[bp_readys__T_218_addr] <= bp_readys__T_218_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_220_en & bp_readys__T_220_mask) begin
      bp_readys[bp_readys__T_220_addr] <= bp_readys__T_220_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_222_en & bp_readys__T_222_mask) begin
      bp_readys[bp_readys__T_222_addr] <= bp_readys__T_222_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_224_en & bp_readys__T_224_mask) begin
      bp_readys[bp_readys__T_224_addr] <= bp_readys__T_224_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_226_en & bp_readys__T_226_mask) begin
      bp_readys[bp_readys__T_226_addr] <= bp_readys__T_226_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_228_en & bp_readys__T_228_mask) begin
      bp_readys[bp_readys__T_228_addr] <= bp_readys__T_228_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_230_en & bp_readys__T_230_mask) begin
      bp_readys[bp_readys__T_230_addr] <= bp_readys__T_230_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_232_en & bp_readys__T_232_mask) begin
      bp_readys[bp_readys__T_232_addr] <= bp_readys__T_232_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_234_en & bp_readys__T_234_mask) begin
      bp_readys[bp_readys__T_234_addr] <= bp_readys__T_234_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_236_en & bp_readys__T_236_mask) begin
      bp_readys[bp_readys__T_236_addr] <= bp_readys__T_236_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_238_en & bp_readys__T_238_mask) begin
      bp_readys[bp_readys__T_238_addr] <= bp_readys__T_238_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_240_en & bp_readys__T_240_mask) begin
      bp_readys[bp_readys__T_240_addr] <= bp_readys__T_240_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_242_en & bp_readys__T_242_mask) begin
      bp_readys[bp_readys__T_242_addr] <= bp_readys__T_242_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_244_en & bp_readys__T_244_mask) begin
      bp_readys[bp_readys__T_244_addr] <= bp_readys__T_244_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_246_en & bp_readys__T_246_mask) begin
      bp_readys[bp_readys__T_246_addr] <= bp_readys__T_246_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_248_en & bp_readys__T_248_mask) begin
      bp_readys[bp_readys__T_248_addr] <= bp_readys__T_248_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_250_en & bp_readys__T_250_mask) begin
      bp_readys[bp_readys__T_250_addr] <= bp_readys__T_250_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_252_en & bp_readys__T_252_mask) begin
      bp_readys[bp_readys__T_252_addr] <= bp_readys__T_252_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_254_en & bp_readys__T_254_mask) begin
      bp_readys[bp_readys__T_254_addr] <= bp_readys__T_254_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_256_en & bp_readys__T_256_mask) begin
      bp_readys[bp_readys__T_256_addr] <= bp_readys__T_256_data; // @[rf.scala 25:22]
    end
    if(bp_readys__T_258_en & bp_readys__T_258_mask) begin
      bp_readys[bp_readys__T_258_addr] <= bp_readys__T_258_data; // @[rf.scala 25:22]
    end
  end
endmodule
module IMemPipe(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [4:0]  io_enq_bits_ex_et,
  input  [4:0]  io_enq_bits_ex_code,
  input  [31:0] io_enq_bits_ex_addr,
  input  [7:0]  io_enq_bits_ex_asid,
  input  [31:0] io_enq_bits_pc,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits_valid,
  output [4:0]  io_deq_bits_bits_ex_et,
  output [4:0]  io_deq_bits_bits_ex_code,
  output [31:0] io_deq_bits_bits_ex_addr,
  output [7:0]  io_deq_bits_bits_ex_asid,
  output [31:0] io_deq_bits_bits_pc,
  input         io_br_flush_valid,
  input         io_ex_flush_valid
);
  reg  queue_valid [0:1]; // @[ifu.scala 26:18]
  reg [31:0] _RAND_0;
  wire  queue_valid__T_21_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_21_addr; // @[ifu.scala 26:18]
  wire  queue_valid_q_head_data; // @[ifu.scala 26:18]
  wire  queue_valid_q_head_addr; // @[ifu.scala 26:18]
  wire  queue_valid_q_head_mask; // @[ifu.scala 26:18]
  wire  queue_valid_q_head_en; // @[ifu.scala 26:18]
  wire  queue_valid__T_12_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_12_addr; // @[ifu.scala 26:18]
  wire  queue_valid__T_12_mask; // @[ifu.scala 26:18]
  wire  queue_valid__T_12_en; // @[ifu.scala 26:18]
  wire  queue_valid__T_15_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_15_addr; // @[ifu.scala 26:18]
  wire  queue_valid__T_15_mask; // @[ifu.scala 26:18]
  wire  queue_valid__T_15_en; // @[ifu.scala 26:18]
  wire  queue_valid__T_25_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_25_addr; // @[ifu.scala 26:18]
  wire  queue_valid__T_25_mask; // @[ifu.scala 26:18]
  wire  queue_valid__T_25_en; // @[ifu.scala 26:18]
  wire  queue_valid__T_26_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_26_addr; // @[ifu.scala 26:18]
  wire  queue_valid__T_26_mask; // @[ifu.scala 26:18]
  wire  queue_valid__T_26_en; // @[ifu.scala 26:18]
  wire  queue_valid__T_31_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_31_addr; // @[ifu.scala 26:18]
  wire  queue_valid__T_31_mask; // @[ifu.scala 26:18]
  wire  queue_valid__T_31_en; // @[ifu.scala 26:18]
  wire  queue_valid__T_33_data; // @[ifu.scala 26:18]
  wire  queue_valid__T_33_addr; // @[ifu.scala 26:18]
  wire  queue_valid__T_33_mask; // @[ifu.scala 26:18]
  wire  queue_valid__T_33_en; // @[ifu.scala 26:18]
  reg [4:0] queue_bits_ex_et [0:1]; // @[ifu.scala 26:18]
  reg [31:0] _RAND_1;
  wire [4:0] queue_bits_ex_et__T_21_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_21_addr; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et_q_head_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et_q_head_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et_q_head_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et_q_head_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et__T_12_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_12_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_12_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_12_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et__T_15_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_15_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_15_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_15_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et__T_25_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_25_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_25_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_25_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et__T_26_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_26_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_26_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_26_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et__T_31_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_31_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_31_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_31_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_et__T_33_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_33_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_33_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_et__T_33_en; // @[ifu.scala 26:18]
  reg [4:0] queue_bits_ex_code [0:1]; // @[ifu.scala 26:18]
  reg [31:0] _RAND_2;
  wire [4:0] queue_bits_ex_code__T_21_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_21_addr; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code_q_head_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code_q_head_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code_q_head_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code_q_head_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code__T_12_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_12_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_12_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_12_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code__T_15_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_15_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_15_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_15_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code__T_25_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_25_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_25_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_25_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code__T_26_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_26_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_26_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_26_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code__T_31_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_31_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_31_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_31_en; // @[ifu.scala 26:18]
  wire [4:0] queue_bits_ex_code__T_33_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_33_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_33_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_code__T_33_en; // @[ifu.scala 26:18]
  reg [31:0] queue_bits_ex_addr [0:1]; // @[ifu.scala 26:18]
  reg [31:0] _RAND_3;
  wire [31:0] queue_bits_ex_addr__T_21_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_21_addr; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr_q_head_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr_q_head_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr_q_head_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr_q_head_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr__T_12_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_12_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_12_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_12_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr__T_15_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_15_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_15_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_15_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr__T_25_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_25_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_25_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_25_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr__T_26_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_26_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_26_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_26_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr__T_31_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_31_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_31_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_31_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_ex_addr__T_33_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_33_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_33_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_addr__T_33_en; // @[ifu.scala 26:18]
  reg [7:0] queue_bits_ex_asid [0:1]; // @[ifu.scala 26:18]
  reg [31:0] _RAND_4;
  wire [7:0] queue_bits_ex_asid__T_21_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_21_addr; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid_q_head_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid_q_head_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid_q_head_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid_q_head_en; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid__T_12_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_12_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_12_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_12_en; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid__T_15_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_15_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_15_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_15_en; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid__T_25_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_25_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_25_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_25_en; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid__T_26_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_26_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_26_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_26_en; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid__T_31_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_31_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_31_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_31_en; // @[ifu.scala 26:18]
  wire [7:0] queue_bits_ex_asid__T_33_data; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_33_addr; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_33_mask; // @[ifu.scala 26:18]
  wire  queue_bits_ex_asid__T_33_en; // @[ifu.scala 26:18]
  reg [31:0] queue_bits_pc [0:1]; // @[ifu.scala 26:18]
  reg [31:0] _RAND_5;
  wire [31:0] queue_bits_pc__T_21_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_21_addr; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc_q_head_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc_q_head_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc_q_head_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc_q_head_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc__T_12_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_12_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_12_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_12_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc__T_15_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_15_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_15_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_15_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc__T_25_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_25_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_25_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_25_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc__T_26_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_26_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_26_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_26_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc__T_31_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_31_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_31_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_31_en; // @[ifu.scala 26:18]
  wire [31:0] queue_bits_pc__T_33_data; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_33_addr; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_33_mask; // @[ifu.scala 26:18]
  wire  queue_bits_pc__T_33_en; // @[ifu.scala 26:18]
  reg  head; // @[ifu.scala 22:21]
  reg [31:0] _RAND_6;
  reg  tail; // @[ifu.scala 23:21]
  reg [31:0] _RAND_7;
  reg  is_full; // @[ifu.scala 24:24]
  reg [31:0] _RAND_8;
  reg  is_empty; // @[ifu.scala 25:25]
  reg [31:0] _RAND_9;
  wire  _T_1 = head + 1'h1; // @[ifu.scala 27:28]
  wire [1:0] _GEN_82 = {{1'd0}, _T_1}; // @[ifu.scala 27:34]
  wire  _T_2 = _GEN_82 == 2'h2; // @[ifu.scala 27:34]
  wire  next_head = _T_2 ? 1'h0 : _T_1; // @[ifu.scala 27:25]
  wire  _T_6 = tail + 1'h1; // @[ifu.scala 27:28]
  wire [1:0] _GEN_83 = {{1'd0}, _T_6}; // @[ifu.scala 27:34]
  wire  _T_7 = _GEN_83 == 2'h2; // @[ifu.scala 27:34]
  wire  next_tail = _T_7 ? 1'h0 : _T_6; // @[ifu.scala 27:25]
  wire  _T_10 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_18 = ~is_full; // @[ifu.scala 39:19]
  wire  _T_20 = ~is_empty; // @[ifu.scala 40:19]
  wire  _T_23 = io_br_flush_valid & _T_10; // @[ifu.scala 50:49]
  wire  _T_24 = io_ex_flush_valid | _T_23; // @[ifu.scala 50:27]
  wire  _T_28 = ~_T_10; // @[ifu.scala 56:36]
  wire  _T_29 = io_br_flush_valid & _T_28; // @[ifu.scala 56:33]
  wire  _T_32 = ~tail; // @[ifu.scala 58:17]
  wire  _T_34 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_35 = next_head == tail; // @[ifu.scala 69:23]
  wire  _T_38 = _T_35 & _T_28; // @[ifu.scala 69:32]
  wire  _GEN_24 = _T_38 | is_full; // @[ifu.scala 69:51]
  wire  _GEN_33 = _T_34 ? 1'h0 : is_empty; // @[ifu.scala 64:26]
  wire  _T_41 = is_full & _T_34; // @[ifu.scala 76:23]
  wire  _T_42 = ~_T_41; // @[ifu.scala 76:13]
  wire  _T_43 = next_tail == head; // @[ifu.scala 77:23]
  wire  _T_45 = ~_T_34; // @[ifu.scala 77:35]
  wire  _T_46 = _T_43 & _T_45; // @[ifu.scala 77:32]
  wire  _GEN_36 = _T_46 | _GEN_33; // @[ifu.scala 77:51]
  wire  _GEN_39 = _T_10 ? _GEN_36 : _GEN_33; // @[ifu.scala 74:26]
  wire  _GEN_42 = _T_29 & tail; // @[ifu.scala 56:52]
  wire  _GEN_46 = _T_29 & _T_32; // @[ifu.scala 56:52]
  wire  _GEN_50 = _T_29 ? 1'h0 : _GEN_39; // @[ifu.scala 56:52]
  wire  _GEN_52 = _T_29 ? 1'h0 : _T_34; // @[ifu.scala 56:52]
  wire  _GEN_62 = _T_24 | _GEN_50; // @[ifu.scala 50:68]
  wire  _T_49 = _T_18 | _T_20; // @[ifu.scala 96:20]
  wire  _T_51 = _T_49 | reset; // @[ifu.scala 96:10]
  wire  _T_52 = ~_T_51; // @[ifu.scala 96:10]
  assign queue_valid__T_21_addr = tail;
  assign queue_valid__T_21_data = queue_valid[queue_valid__T_21_addr]; // @[ifu.scala 26:18]
  assign queue_valid_q_head_data = 1'h1;
  assign queue_valid_q_head_addr = head;
  assign queue_valid_q_head_mask = _T_24 ? 1'h0 : _GEN_52;
  assign queue_valid_q_head_en = 1'h1;
  assign queue_valid__T_12_data = 1'h0;
  assign queue_valid__T_12_addr = 1'h0;
  assign queue_valid__T_12_mask = 1'h1;
  assign queue_valid__T_12_en = reset;
  assign queue_valid__T_15_data = 1'h0;
  assign queue_valid__T_15_addr = 1'h1;
  assign queue_valid__T_15_mask = 1'h1;
  assign queue_valid__T_15_en = reset;
  assign queue_valid__T_25_data = 1'h0;
  assign queue_valid__T_25_addr = 1'h0;
  assign queue_valid__T_25_mask = 1'h1;
  assign queue_valid__T_25_en = io_ex_flush_valid | _T_23;
  assign queue_valid__T_26_data = 1'h0;
  assign queue_valid__T_26_addr = 1'h1;
  assign queue_valid__T_26_mask = 1'h1;
  assign queue_valid__T_26_en = io_ex_flush_valid | _T_23;
  assign queue_valid__T_31_data = 1'h0;
  assign queue_valid__T_31_addr = 1'h0;
  assign queue_valid__T_31_mask = 1'h1;
  assign queue_valid__T_31_en = _T_24 ? 1'h0 : _GEN_42;
  assign queue_valid__T_33_data = 1'h0;
  assign queue_valid__T_33_addr = 1'h1;
  assign queue_valid__T_33_mask = 1'h1;
  assign queue_valid__T_33_en = _T_24 ? 1'h0 : _GEN_46;
  assign queue_bits_ex_et__T_21_addr = tail;
  assign queue_bits_ex_et__T_21_data = queue_bits_ex_et[queue_bits_ex_et__T_21_addr]; // @[ifu.scala 26:18]
  assign queue_bits_ex_et_q_head_data = io_enq_bits_ex_et;
  assign queue_bits_ex_et_q_head_addr = head;
  assign queue_bits_ex_et_q_head_mask = _T_24 ? 1'h0 : _GEN_52;
  assign queue_bits_ex_et_q_head_en = 1'h1;
  assign queue_bits_ex_et__T_12_data = 5'h0;
  assign queue_bits_ex_et__T_12_addr = 1'h0;
  assign queue_bits_ex_et__T_12_mask = 1'h1;
  assign queue_bits_ex_et__T_12_en = reset;
  assign queue_bits_ex_et__T_15_data = 5'h0;
  assign queue_bits_ex_et__T_15_addr = 1'h1;
  assign queue_bits_ex_et__T_15_mask = 1'h1;
  assign queue_bits_ex_et__T_15_en = reset;
  assign queue_bits_ex_et__T_25_data = 5'h0;
  assign queue_bits_ex_et__T_25_addr = 1'h0;
  assign queue_bits_ex_et__T_25_mask = 1'h0;
  assign queue_bits_ex_et__T_25_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_et__T_26_data = 5'h0;
  assign queue_bits_ex_et__T_26_addr = 1'h1;
  assign queue_bits_ex_et__T_26_mask = 1'h0;
  assign queue_bits_ex_et__T_26_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_et__T_31_data = 5'h0;
  assign queue_bits_ex_et__T_31_addr = 1'h0;
  assign queue_bits_ex_et__T_31_mask = 1'h0;
  assign queue_bits_ex_et__T_31_en = _T_24 ? 1'h0 : _GEN_42;
  assign queue_bits_ex_et__T_33_data = 5'h0;
  assign queue_bits_ex_et__T_33_addr = 1'h1;
  assign queue_bits_ex_et__T_33_mask = 1'h0;
  assign queue_bits_ex_et__T_33_en = _T_24 ? 1'h0 : _GEN_46;
  assign queue_bits_ex_code__T_21_addr = tail;
  assign queue_bits_ex_code__T_21_data = queue_bits_ex_code[queue_bits_ex_code__T_21_addr]; // @[ifu.scala 26:18]
  assign queue_bits_ex_code_q_head_data = io_enq_bits_ex_code;
  assign queue_bits_ex_code_q_head_addr = head;
  assign queue_bits_ex_code_q_head_mask = _T_24 ? 1'h0 : _GEN_52;
  assign queue_bits_ex_code_q_head_en = 1'h1;
  assign queue_bits_ex_code__T_12_data = 5'h0;
  assign queue_bits_ex_code__T_12_addr = 1'h0;
  assign queue_bits_ex_code__T_12_mask = 1'h1;
  assign queue_bits_ex_code__T_12_en = reset;
  assign queue_bits_ex_code__T_15_data = 5'h0;
  assign queue_bits_ex_code__T_15_addr = 1'h1;
  assign queue_bits_ex_code__T_15_mask = 1'h1;
  assign queue_bits_ex_code__T_15_en = reset;
  assign queue_bits_ex_code__T_25_data = 5'h0;
  assign queue_bits_ex_code__T_25_addr = 1'h0;
  assign queue_bits_ex_code__T_25_mask = 1'h0;
  assign queue_bits_ex_code__T_25_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_code__T_26_data = 5'h0;
  assign queue_bits_ex_code__T_26_addr = 1'h1;
  assign queue_bits_ex_code__T_26_mask = 1'h0;
  assign queue_bits_ex_code__T_26_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_code__T_31_data = 5'h0;
  assign queue_bits_ex_code__T_31_addr = 1'h0;
  assign queue_bits_ex_code__T_31_mask = 1'h0;
  assign queue_bits_ex_code__T_31_en = _T_24 ? 1'h0 : _GEN_42;
  assign queue_bits_ex_code__T_33_data = 5'h0;
  assign queue_bits_ex_code__T_33_addr = 1'h1;
  assign queue_bits_ex_code__T_33_mask = 1'h0;
  assign queue_bits_ex_code__T_33_en = _T_24 ? 1'h0 : _GEN_46;
  assign queue_bits_ex_addr__T_21_addr = tail;
  assign queue_bits_ex_addr__T_21_data = queue_bits_ex_addr[queue_bits_ex_addr__T_21_addr]; // @[ifu.scala 26:18]
  assign queue_bits_ex_addr_q_head_data = io_enq_bits_ex_addr;
  assign queue_bits_ex_addr_q_head_addr = head;
  assign queue_bits_ex_addr_q_head_mask = _T_24 ? 1'h0 : _GEN_52;
  assign queue_bits_ex_addr_q_head_en = 1'h1;
  assign queue_bits_ex_addr__T_12_data = 32'h0;
  assign queue_bits_ex_addr__T_12_addr = 1'h0;
  assign queue_bits_ex_addr__T_12_mask = 1'h1;
  assign queue_bits_ex_addr__T_12_en = reset;
  assign queue_bits_ex_addr__T_15_data = 32'h0;
  assign queue_bits_ex_addr__T_15_addr = 1'h1;
  assign queue_bits_ex_addr__T_15_mask = 1'h1;
  assign queue_bits_ex_addr__T_15_en = reset;
  assign queue_bits_ex_addr__T_25_data = 32'h0;
  assign queue_bits_ex_addr__T_25_addr = 1'h0;
  assign queue_bits_ex_addr__T_25_mask = 1'h0;
  assign queue_bits_ex_addr__T_25_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_addr__T_26_data = 32'h0;
  assign queue_bits_ex_addr__T_26_addr = 1'h1;
  assign queue_bits_ex_addr__T_26_mask = 1'h0;
  assign queue_bits_ex_addr__T_26_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_addr__T_31_data = 32'h0;
  assign queue_bits_ex_addr__T_31_addr = 1'h0;
  assign queue_bits_ex_addr__T_31_mask = 1'h0;
  assign queue_bits_ex_addr__T_31_en = _T_24 ? 1'h0 : _GEN_42;
  assign queue_bits_ex_addr__T_33_data = 32'h0;
  assign queue_bits_ex_addr__T_33_addr = 1'h1;
  assign queue_bits_ex_addr__T_33_mask = 1'h0;
  assign queue_bits_ex_addr__T_33_en = _T_24 ? 1'h0 : _GEN_46;
  assign queue_bits_ex_asid__T_21_addr = tail;
  assign queue_bits_ex_asid__T_21_data = queue_bits_ex_asid[queue_bits_ex_asid__T_21_addr]; // @[ifu.scala 26:18]
  assign queue_bits_ex_asid_q_head_data = io_enq_bits_ex_asid;
  assign queue_bits_ex_asid_q_head_addr = head;
  assign queue_bits_ex_asid_q_head_mask = _T_24 ? 1'h0 : _GEN_52;
  assign queue_bits_ex_asid_q_head_en = 1'h1;
  assign queue_bits_ex_asid__T_12_data = 8'h0;
  assign queue_bits_ex_asid__T_12_addr = 1'h0;
  assign queue_bits_ex_asid__T_12_mask = 1'h1;
  assign queue_bits_ex_asid__T_12_en = reset;
  assign queue_bits_ex_asid__T_15_data = 8'h0;
  assign queue_bits_ex_asid__T_15_addr = 1'h1;
  assign queue_bits_ex_asid__T_15_mask = 1'h1;
  assign queue_bits_ex_asid__T_15_en = reset;
  assign queue_bits_ex_asid__T_25_data = 8'h0;
  assign queue_bits_ex_asid__T_25_addr = 1'h0;
  assign queue_bits_ex_asid__T_25_mask = 1'h0;
  assign queue_bits_ex_asid__T_25_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_asid__T_26_data = 8'h0;
  assign queue_bits_ex_asid__T_26_addr = 1'h1;
  assign queue_bits_ex_asid__T_26_mask = 1'h0;
  assign queue_bits_ex_asid__T_26_en = io_ex_flush_valid | _T_23;
  assign queue_bits_ex_asid__T_31_data = 8'h0;
  assign queue_bits_ex_asid__T_31_addr = 1'h0;
  assign queue_bits_ex_asid__T_31_mask = 1'h0;
  assign queue_bits_ex_asid__T_31_en = _T_24 ? 1'h0 : _GEN_42;
  assign queue_bits_ex_asid__T_33_data = 8'h0;
  assign queue_bits_ex_asid__T_33_addr = 1'h1;
  assign queue_bits_ex_asid__T_33_mask = 1'h0;
  assign queue_bits_ex_asid__T_33_en = _T_24 ? 1'h0 : _GEN_46;
  assign queue_bits_pc__T_21_addr = tail;
  assign queue_bits_pc__T_21_data = queue_bits_pc[queue_bits_pc__T_21_addr]; // @[ifu.scala 26:18]
  assign queue_bits_pc_q_head_data = io_enq_bits_pc;
  assign queue_bits_pc_q_head_addr = head;
  assign queue_bits_pc_q_head_mask = _T_24 ? 1'h0 : _GEN_52;
  assign queue_bits_pc_q_head_en = 1'h1;
  assign queue_bits_pc__T_12_data = 32'h0;
  assign queue_bits_pc__T_12_addr = 1'h0;
  assign queue_bits_pc__T_12_mask = 1'h1;
  assign queue_bits_pc__T_12_en = reset;
  assign queue_bits_pc__T_15_data = 32'h0;
  assign queue_bits_pc__T_15_addr = 1'h1;
  assign queue_bits_pc__T_15_mask = 1'h1;
  assign queue_bits_pc__T_15_en = reset;
  assign queue_bits_pc__T_25_data = 32'h0;
  assign queue_bits_pc__T_25_addr = 1'h0;
  assign queue_bits_pc__T_25_mask = 1'h0;
  assign queue_bits_pc__T_25_en = io_ex_flush_valid | _T_23;
  assign queue_bits_pc__T_26_data = 32'h0;
  assign queue_bits_pc__T_26_addr = 1'h1;
  assign queue_bits_pc__T_26_mask = 1'h0;
  assign queue_bits_pc__T_26_en = io_ex_flush_valid | _T_23;
  assign queue_bits_pc__T_31_data = 32'h0;
  assign queue_bits_pc__T_31_addr = 1'h0;
  assign queue_bits_pc__T_31_mask = 1'h0;
  assign queue_bits_pc__T_31_en = _T_24 ? 1'h0 : _GEN_42;
  assign queue_bits_pc__T_33_data = 32'h0;
  assign queue_bits_pc__T_33_addr = 1'h1;
  assign queue_bits_pc__T_33_mask = 1'h0;
  assign queue_bits_pc__T_33_en = _T_24 ? 1'h0 : _GEN_46;
  assign io_enq_ready = _T_18 | io_deq_ready; // @[ifu.scala 39:16]
  assign io_deq_valid = ~is_empty; // @[ifu.scala 40:16]
  assign io_deq_bits_valid = queue_valid__T_21_data; // @[ifu.scala 41:15]
  assign io_deq_bits_bits_ex_et = queue_bits_ex_et__T_21_data; // @[ifu.scala 41:15]
  assign io_deq_bits_bits_ex_code = queue_bits_ex_code__T_21_data; // @[ifu.scala 41:15]
  assign io_deq_bits_bits_ex_addr = queue_bits_ex_addr__T_21_data; // @[ifu.scala 41:15]
  assign io_deq_bits_bits_ex_asid = queue_bits_ex_asid__T_21_data; // @[ifu.scala 41:15]
  assign io_deq_bits_bits_pc = queue_bits_pc__T_21_data; // @[ifu.scala 41:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    queue_valid[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    queue_bits_ex_et[initvar] = _RAND_1[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    queue_bits_ex_code[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    queue_bits_ex_addr[initvar] = _RAND_3[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    queue_bits_ex_asid[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    queue_bits_pc[initvar] = _RAND_5[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  head = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tail = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  is_full = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  is_empty = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(queue_valid_q_head_en & queue_valid_q_head_mask) begin
      queue_valid[queue_valid_q_head_addr] <= queue_valid_q_head_data; // @[ifu.scala 26:18]
    end
    if(queue_valid__T_12_en & queue_valid__T_12_mask) begin
      queue_valid[queue_valid__T_12_addr] <= queue_valid__T_12_data; // @[ifu.scala 26:18]
    end
    if(queue_valid__T_15_en & queue_valid__T_15_mask) begin
      queue_valid[queue_valid__T_15_addr] <= queue_valid__T_15_data; // @[ifu.scala 26:18]
    end
    if(queue_valid__T_25_en & queue_valid__T_25_mask) begin
      queue_valid[queue_valid__T_25_addr] <= queue_valid__T_25_data; // @[ifu.scala 26:18]
    end
    if(queue_valid__T_26_en & queue_valid__T_26_mask) begin
      queue_valid[queue_valid__T_26_addr] <= queue_valid__T_26_data; // @[ifu.scala 26:18]
    end
    if(queue_valid__T_31_en & queue_valid__T_31_mask) begin
      queue_valid[queue_valid__T_31_addr] <= queue_valid__T_31_data; // @[ifu.scala 26:18]
    end
    if(queue_valid__T_33_en & queue_valid__T_33_mask) begin
      queue_valid[queue_valid__T_33_addr] <= queue_valid__T_33_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et_q_head_en & queue_bits_ex_et_q_head_mask) begin
      queue_bits_ex_et[queue_bits_ex_et_q_head_addr] <= queue_bits_ex_et_q_head_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et__T_12_en & queue_bits_ex_et__T_12_mask) begin
      queue_bits_ex_et[queue_bits_ex_et__T_12_addr] <= queue_bits_ex_et__T_12_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et__T_15_en & queue_bits_ex_et__T_15_mask) begin
      queue_bits_ex_et[queue_bits_ex_et__T_15_addr] <= queue_bits_ex_et__T_15_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et__T_25_en & queue_bits_ex_et__T_25_mask) begin
      queue_bits_ex_et[queue_bits_ex_et__T_25_addr] <= queue_bits_ex_et__T_25_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et__T_26_en & queue_bits_ex_et__T_26_mask) begin
      queue_bits_ex_et[queue_bits_ex_et__T_26_addr] <= queue_bits_ex_et__T_26_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et__T_31_en & queue_bits_ex_et__T_31_mask) begin
      queue_bits_ex_et[queue_bits_ex_et__T_31_addr] <= queue_bits_ex_et__T_31_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_et__T_33_en & queue_bits_ex_et__T_33_mask) begin
      queue_bits_ex_et[queue_bits_ex_et__T_33_addr] <= queue_bits_ex_et__T_33_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code_q_head_en & queue_bits_ex_code_q_head_mask) begin
      queue_bits_ex_code[queue_bits_ex_code_q_head_addr] <= queue_bits_ex_code_q_head_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code__T_12_en & queue_bits_ex_code__T_12_mask) begin
      queue_bits_ex_code[queue_bits_ex_code__T_12_addr] <= queue_bits_ex_code__T_12_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code__T_15_en & queue_bits_ex_code__T_15_mask) begin
      queue_bits_ex_code[queue_bits_ex_code__T_15_addr] <= queue_bits_ex_code__T_15_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code__T_25_en & queue_bits_ex_code__T_25_mask) begin
      queue_bits_ex_code[queue_bits_ex_code__T_25_addr] <= queue_bits_ex_code__T_25_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code__T_26_en & queue_bits_ex_code__T_26_mask) begin
      queue_bits_ex_code[queue_bits_ex_code__T_26_addr] <= queue_bits_ex_code__T_26_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code__T_31_en & queue_bits_ex_code__T_31_mask) begin
      queue_bits_ex_code[queue_bits_ex_code__T_31_addr] <= queue_bits_ex_code__T_31_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_code__T_33_en & queue_bits_ex_code__T_33_mask) begin
      queue_bits_ex_code[queue_bits_ex_code__T_33_addr] <= queue_bits_ex_code__T_33_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr_q_head_en & queue_bits_ex_addr_q_head_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr_q_head_addr] <= queue_bits_ex_addr_q_head_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr__T_12_en & queue_bits_ex_addr__T_12_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr__T_12_addr] <= queue_bits_ex_addr__T_12_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr__T_15_en & queue_bits_ex_addr__T_15_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr__T_15_addr] <= queue_bits_ex_addr__T_15_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr__T_25_en & queue_bits_ex_addr__T_25_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr__T_25_addr] <= queue_bits_ex_addr__T_25_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr__T_26_en & queue_bits_ex_addr__T_26_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr__T_26_addr] <= queue_bits_ex_addr__T_26_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr__T_31_en & queue_bits_ex_addr__T_31_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr__T_31_addr] <= queue_bits_ex_addr__T_31_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_addr__T_33_en & queue_bits_ex_addr__T_33_mask) begin
      queue_bits_ex_addr[queue_bits_ex_addr__T_33_addr] <= queue_bits_ex_addr__T_33_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid_q_head_en & queue_bits_ex_asid_q_head_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid_q_head_addr] <= queue_bits_ex_asid_q_head_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid__T_12_en & queue_bits_ex_asid__T_12_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid__T_12_addr] <= queue_bits_ex_asid__T_12_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid__T_15_en & queue_bits_ex_asid__T_15_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid__T_15_addr] <= queue_bits_ex_asid__T_15_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid__T_25_en & queue_bits_ex_asid__T_25_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid__T_25_addr] <= queue_bits_ex_asid__T_25_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid__T_26_en & queue_bits_ex_asid__T_26_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid__T_26_addr] <= queue_bits_ex_asid__T_26_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid__T_31_en & queue_bits_ex_asid__T_31_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid__T_31_addr] <= queue_bits_ex_asid__T_31_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_ex_asid__T_33_en & queue_bits_ex_asid__T_33_mask) begin
      queue_bits_ex_asid[queue_bits_ex_asid__T_33_addr] <= queue_bits_ex_asid__T_33_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc_q_head_en & queue_bits_pc_q_head_mask) begin
      queue_bits_pc[queue_bits_pc_q_head_addr] <= queue_bits_pc_q_head_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc__T_12_en & queue_bits_pc__T_12_mask) begin
      queue_bits_pc[queue_bits_pc__T_12_addr] <= queue_bits_pc__T_12_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc__T_15_en & queue_bits_pc__T_15_mask) begin
      queue_bits_pc[queue_bits_pc__T_15_addr] <= queue_bits_pc__T_15_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc__T_25_en & queue_bits_pc__T_25_mask) begin
      queue_bits_pc[queue_bits_pc__T_25_addr] <= queue_bits_pc__T_25_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc__T_26_en & queue_bits_pc__T_26_mask) begin
      queue_bits_pc[queue_bits_pc__T_26_addr] <= queue_bits_pc__T_26_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc__T_31_en & queue_bits_pc__T_31_mask) begin
      queue_bits_pc[queue_bits_pc__T_31_addr] <= queue_bits_pc__T_31_data; // @[ifu.scala 26:18]
    end
    if(queue_bits_pc__T_33_en & queue_bits_pc__T_33_mask) begin
      queue_bits_pc[queue_bits_pc__T_33_addr] <= queue_bits_pc__T_33_data; // @[ifu.scala 26:18]
    end
    if (reset) begin
      head <= 1'h0;
    end else if (_T_24) begin
      head <= 1'h0;
    end else if (_T_29) begin
      if (_T_7) begin
        head <= 1'h0;
      end else begin
        head <= _T_6;
      end
    end else if (_T_34) begin
      if (_T_2) begin
        head <= 1'h0;
      end else begin
        head <= _T_1;
      end
    end
    if (reset) begin
      tail <= 1'h0;
    end else if (_T_24) begin
      tail <= 1'h0;
    end else if (!(_T_29)) begin
      if (_T_10) begin
        if (_T_7) begin
          tail <= 1'h0;
        end else begin
          tail <= _T_6;
        end
      end
    end
    if (reset) begin
      is_full <= 1'h0;
    end else if (_T_24) begin
      is_full <= 1'h0;
    end else if (_T_29) begin
      is_full <= 1'h0;
    end else if (_T_10) begin
      if (_T_42) begin
        is_full <= 1'h0;
      end else if (_T_34) begin
        is_full <= _GEN_24;
      end
    end else if (_T_34) begin
      is_full <= _GEN_24;
    end
    is_empty <= reset | _GEN_62;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_52) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ifu.scala:96 assert (!is_full || !is_empty)\n"); // @[ifu.scala 96:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_52) begin
          $fatal; // @[ifu.scala 96:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module IFU(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output        io_imem_req_bits_is_cached,
  output [31:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [31:0] io_imem_resp_bits_data,
  input         io_iaddr_req_ready,
  output        io_iaddr_req_valid,
  output [31:0] io_iaddr_req_bits_vaddr,
  output        io_iaddr_resp_ready,
  input         io_iaddr_resp_valid,
  input  [31:0] io_iaddr_resp_bits_paddr,
  input         io_iaddr_resp_bits_is_cached,
  input  [4:0]  io_iaddr_resp_bits_ex_et,
  input  [4:0]  io_iaddr_resp_bits_ex_code,
  input  [31:0] io_iaddr_resp_bits_ex_addr,
  input  [7:0]  io_iaddr_resp_bits_ex_asid,
  input         io_fu_out_ready,
  output        io_fu_out_valid,
  output [31:0] io_fu_out_bits_pc,
  output [31:0] io_fu_out_bits_instr,
  output [4:0]  io_fu_out_bits_ex_et,
  output [4:0]  io_fu_out_bits_ex_code,
  output [31:0] io_fu_out_bits_ex_addr,
  output [7:0]  io_fu_out_bits_ex_asid,
  input         io_br_flush_valid,
  input  [31:0] io_br_flush_bits_br_target,
  input         io_ex_flush_valid,
  input  [31:0] io_ex_flush_bits_br_target
);
  wire  s1_datas_clock; // @[ifu.scala 141:24]
  wire  s1_datas_reset; // @[ifu.scala 141:24]
  wire  s1_datas_io_enq_ready; // @[ifu.scala 141:24]
  wire  s1_datas_io_enq_valid; // @[ifu.scala 141:24]
  wire [4:0] s1_datas_io_enq_bits_ex_et; // @[ifu.scala 141:24]
  wire [4:0] s1_datas_io_enq_bits_ex_code; // @[ifu.scala 141:24]
  wire [31:0] s1_datas_io_enq_bits_ex_addr; // @[ifu.scala 141:24]
  wire [7:0] s1_datas_io_enq_bits_ex_asid; // @[ifu.scala 141:24]
  wire [31:0] s1_datas_io_enq_bits_pc; // @[ifu.scala 141:24]
  wire  s1_datas_io_deq_ready; // @[ifu.scala 141:24]
  wire  s1_datas_io_deq_valid; // @[ifu.scala 141:24]
  wire  s1_datas_io_deq_bits_valid; // @[ifu.scala 141:24]
  wire [4:0] s1_datas_io_deq_bits_bits_ex_et; // @[ifu.scala 141:24]
  wire [4:0] s1_datas_io_deq_bits_bits_ex_code; // @[ifu.scala 141:24]
  wire [31:0] s1_datas_io_deq_bits_bits_ex_addr; // @[ifu.scala 141:24]
  wire [7:0] s1_datas_io_deq_bits_bits_ex_asid; // @[ifu.scala 141:24]
  wire [31:0] s1_datas_io_deq_bits_bits_pc; // @[ifu.scala 141:24]
  wire  s1_datas_io_br_flush_valid; // @[ifu.scala 141:24]
  wire  s1_datas_io_ex_flush_valid; // @[ifu.scala 141:24]
  reg [31:0] pc; // @[ifu.scala 115:19]
  reg [31:0] _RAND_0;
  wire  pc_misaligned = pc[1:0] != 2'h0; // @[ifu.scala 116:32]
  reg  s0_bad_if; // @[ifu.scala 117:26]
  reg [31:0] _RAND_1;
  wire  _T_1 = io_iaddr_req_ready & io_iaddr_req_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _T_3 = pc + 32'h4; // @[ifu.scala 121:32]
  wire  _T_9 = io_iaddr_req_valid & pc_misaligned; // @[ifu.scala 124:35]
  wire  _GEN_0 = _T_9 | s0_bad_if; // @[ifu.scala 124:56]
  wire  _T_10 = ~io_ex_flush_valid; // @[ifu.scala 129:30]
  wire  _T_12 = ~io_br_flush_valid; // @[ifu.scala 129:52]
  wire  _T_13 = _T_10 & _T_12; // @[ifu.scala 129:49]
  wire  _T_14 = ~s0_bad_if; // @[ifu.scala 129:74]
  reg [31:0] s1_in_pc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  wire  _T_20 = io_iaddr_resp_bits_ex_et != 5'h0; // @[ifu.scala 143:53]
  wire  s1_ex_in = io_iaddr_resp_valid & _T_20; // @[ifu.scala 143:38]
  wire  s1_out_has_ex = s1_datas_io_deq_bits_bits_ex_et != 5'h0; // @[ifu.scala 144:41]
  wire  _T_21 = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_23 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_26 = io_iaddr_resp_valid & _T_10; // @[ifu.scala 151:44]
  wire  _T_27 = io_iaddr_resp_bits_ex_et == 5'h0; // @[ifu.scala 151:81]
  wire  _T_29 = io_imem_resp_valid | s1_out_has_ex; // @[ifu.scala 161:42]
  wire  _T_30 = _T_29 & s1_datas_io_deq_bits_valid; // @[ifu.scala 161:60]
  IMemPipe s1_datas ( // @[ifu.scala 141:24]
    .clock(s1_datas_clock),
    .reset(s1_datas_reset),
    .io_enq_ready(s1_datas_io_enq_ready),
    .io_enq_valid(s1_datas_io_enq_valid),
    .io_enq_bits_ex_et(s1_datas_io_enq_bits_ex_et),
    .io_enq_bits_ex_code(s1_datas_io_enq_bits_ex_code),
    .io_enq_bits_ex_addr(s1_datas_io_enq_bits_ex_addr),
    .io_enq_bits_ex_asid(s1_datas_io_enq_bits_ex_asid),
    .io_enq_bits_pc(s1_datas_io_enq_bits_pc),
    .io_deq_ready(s1_datas_io_deq_ready),
    .io_deq_valid(s1_datas_io_deq_valid),
    .io_deq_bits_valid(s1_datas_io_deq_bits_valid),
    .io_deq_bits_bits_ex_et(s1_datas_io_deq_bits_bits_ex_et),
    .io_deq_bits_bits_ex_code(s1_datas_io_deq_bits_bits_ex_code),
    .io_deq_bits_bits_ex_addr(s1_datas_io_deq_bits_bits_ex_addr),
    .io_deq_bits_bits_ex_asid(s1_datas_io_deq_bits_bits_ex_asid),
    .io_deq_bits_bits_pc(s1_datas_io_deq_bits_bits_pc),
    .io_br_flush_valid(s1_datas_io_br_flush_valid),
    .io_ex_flush_valid(s1_datas_io_ex_flush_valid)
  );
  assign io_imem_req_valid = _T_26 & _T_27; // @[ifu.scala 151:21]
  assign io_imem_req_bits_is_cached = io_iaddr_resp_bits_is_cached; // @[ifu.scala 152:30]
  assign io_imem_req_bits_addr = io_iaddr_resp_bits_paddr; // @[ifu.scala 153:26]
  assign io_imem_resp_ready = io_fu_out_ready; // @[ifu.scala 158:22]
  assign io_iaddr_req_valid = _T_13 & _T_14; // @[ifu.scala 129:22]
  assign io_iaddr_req_bits_vaddr = pc; // @[ifu.scala 133:27]
  assign io_iaddr_resp_ready = io_imem_req_ready; // @[ifu.scala 134:23]
  assign io_fu_out_valid = _T_30 & _T_10; // @[ifu.scala 161:19]
  assign io_fu_out_bits_pc = s1_datas_io_deq_bits_bits_pc; // @[ifu.scala 162:21]
  assign io_fu_out_bits_instr = s1_out_has_ex ? 32'h0 : io_imem_resp_bits_data; // @[ifu.scala 163:24]
  assign io_fu_out_bits_ex_et = s1_datas_io_deq_bits_bits_ex_et; // @[ifu.scala 164:21]
  assign io_fu_out_bits_ex_code = s1_datas_io_deq_bits_bits_ex_code; // @[ifu.scala 164:21]
  assign io_fu_out_bits_ex_addr = s1_datas_io_deq_bits_bits_ex_addr; // @[ifu.scala 164:21]
  assign io_fu_out_bits_ex_asid = s1_datas_io_deq_bits_bits_ex_asid; // @[ifu.scala 164:21]
  assign s1_datas_clock = clock;
  assign s1_datas_reset = reset;
  assign s1_datas_io_enq_valid = _T_21 | s1_ex_in; // @[ifu.scala 145:25]
  assign s1_datas_io_enq_bits_ex_et = io_iaddr_resp_bits_ex_et; // @[ifu.scala 146:24]
  assign s1_datas_io_enq_bits_ex_code = io_iaddr_resp_bits_ex_code; // @[ifu.scala 146:24]
  assign s1_datas_io_enq_bits_ex_addr = io_iaddr_resp_bits_ex_addr; // @[ifu.scala 146:24]
  assign s1_datas_io_enq_bits_ex_asid = io_iaddr_resp_bits_ex_asid; // @[ifu.scala 146:24]
  assign s1_datas_io_enq_bits_pc = s1_in_pc; // @[ifu.scala 146:24]
  assign s1_datas_io_deq_ready = _T_23 | s1_out_has_ex; // @[ifu.scala 147:25]
  assign s1_datas_io_br_flush_valid = io_br_flush_valid; // @[ifu.scala 148:24]
  assign s1_datas_io_ex_flush_valid = io_ex_flush_valid; // @[ifu.scala 149:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  s0_bad_if = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  s1_in_pc = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'hbfc00000;
    end else if (io_ex_flush_valid) begin
      pc <= io_ex_flush_bits_br_target;
    end else if (io_br_flush_valid) begin
      pc <= io_br_flush_bits_br_target;
    end else if (_T_1) begin
      pc <= _T_3;
    end
    if (reset) begin
      s0_bad_if <= 1'h0;
    end else if (io_ex_flush_valid) begin
      s0_bad_if <= 1'h0;
    end else begin
      s0_bad_if <= _GEN_0;
    end
    if (reset) begin
      s1_in_pc <= 32'h0;
    end else if (_T_1) begin
      s1_in_pc <= pc;
    end
  end
endmodule
module BRU(
  input         io_fu_in_valid,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input         io_fu_in_bits_wb_is_ds,
  input  [4:0]  io_fu_in_bits_ops_fu_op,
  input  [31:0] io_fu_in_bits_ops_op1,
  input  [31:0] io_fu_in_bits_ops_op2,
  output        io_fu_out_valid,
  output        io_fu_out_bits_wb_v,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output        io_fu_out_bits_wb_wen,
  output [31:0] io_fu_out_bits_wb_data,
  output        io_fu_out_bits_wb_is_ds,
  output [31:0] io_fu_out_bits_br_target
);
  wire [15:0] _T_1 = {io_fu_in_bits_wb_instr_rd_idx,io_fu_in_bits_wb_instr_shamt,io_fu_in_bits_wb_instr_func}; // @[Cat.scala 29:58]
  wire [15:0] _T_3 = {io_fu_in_bits_wb_instr_rd_idx,io_fu_in_bits_wb_instr_shamt,io_fu_in_bits_wb_instr_func}; // @[bru.scala 19:32]
  wire [31:0] simm = {{16{_T_3[15]}},_T_3}; // @[bru.scala 19:54]
  wire [31:0] _T_5 = io_fu_in_bits_wb_pc + 32'h4; // @[bru.scala 23:16]
  wire [33:0] _T_6 = {simm, 2'h0}; // @[bru.scala 23:30]
  wire [33:0] _GEN_0 = {{2'd0}, _T_5}; // @[bru.scala 23:22]
  wire [33:0] _T_8 = _GEN_0 + _T_6; // @[bru.scala 23:22]
  wire [31:0] Ia = _T_8[31:0]; // @[bru.scala 23:36]
  wire [17:0] _T_19 = {_T_1, 2'h0}; // @[bru.scala 25:42]
  wire [31:0] _T_20 = {{14{_T_19[17]}},_T_19}; // @[bru.scala 25:55]
  wire [31:0] _T_22 = io_fu_in_bits_wb_pc + _T_20; // @[bru.scala 25:15]
  wire [31:0] Za = _T_22 + 32'h4; // @[bru.scala 25:62]
  wire  _T_24 = io_fu_in_bits_ops_op1 == io_fu_in_bits_ops_op2; // @[bru.scala 29:25]
  wire [33:0] _T_26 = {_T_24,1'h0,Ia}; // @[Cat.scala 29:58]
  wire  _T_27 = io_fu_in_bits_ops_op1 != io_fu_in_bits_ops_op2; // @[bru.scala 30:25]
  wire [33:0] _T_29 = {_T_27,1'h0,Ia}; // @[Cat.scala 29:58]
  wire  _T_31 = $signed(io_fu_in_bits_ops_op1) <= 32'sh0; // @[bru.scala 31:32]
  wire [33:0] _T_33 = {_T_31,1'h0,Ia}; // @[Cat.scala 29:58]
  wire  _T_35 = $signed(io_fu_in_bits_ops_op1) >= 32'sh0; // @[bru.scala 32:32]
  wire [33:0] _T_37 = {_T_35,1'h0,Ia}; // @[Cat.scala 29:58]
  wire  _T_39 = $signed(io_fu_in_bits_ops_op1) < 32'sh0; // @[bru.scala 33:32]
  wire [33:0] _T_41 = {_T_39,1'h0,Ia}; // @[Cat.scala 29:58]
  wire  _T_43 = $signed(io_fu_in_bits_ops_op1) > 32'sh0; // @[bru.scala 34:32]
  wire [33:0] _T_45 = {_T_43,1'h0,Ia}; // @[Cat.scala 29:58]
  wire [33:0] _T_49 = {_T_35,1'h1,Za}; // @[Cat.scala 29:58]
  wire [33:0] _T_53 = {_T_39,1'h1,Za}; // @[Cat.scala 29:58]
  wire [34:0] _T_56 = {2'h3,1'h0,io_fu_in_bits_wb_pc[31:28],io_fu_in_bits_wb_instr_rs_idx,io_fu_in_bits_wb_instr_rt_idx,io_fu_in_bits_wb_instr_rd_idx,io_fu_in_bits_wb_instr_shamt,io_fu_in_bits_wb_instr_func,2'h0}; // @[Cat.scala 29:58]
  wire [34:0] _T_59 = {2'h3,1'h1,io_fu_in_bits_wb_pc[31:28],io_fu_in_bits_wb_instr_rs_idx,io_fu_in_bits_wb_instr_rt_idx,io_fu_in_bits_wb_instr_rd_idx,io_fu_in_bits_wb_instr_shamt,io_fu_in_bits_wb_instr_func,2'h0}; // @[Cat.scala 29:58]
  wire [34:0] _T_62 = {2'h3,1'h0,io_fu_in_bits_ops_op1}; // @[Cat.scala 29:58]
  wire [34:0] _T_65 = {2'h3,1'h1,io_fu_in_bits_ops_op1}; // @[Cat.scala 29:58]
  wire  _T_66 = 5'hb == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_67 = _T_66 ? _T_65 : 35'h0; // @[Mux.scala 68:16]
  wire  _T_68 = 5'ha == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_69 = _T_68 ? _T_62 : _T_67; // @[Mux.scala 68:16]
  wire  _T_70 = 5'h9 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_71 = _T_70 ? _T_59 : _T_69; // @[Mux.scala 68:16]
  wire  _T_72 = 5'h8 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_73 = _T_72 ? _T_56 : _T_71; // @[Mux.scala 68:16]
  wire  _T_74 = 5'h7 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_75 = _T_74 ? {{1'd0}, _T_53} : _T_73; // @[Mux.scala 68:16]
  wire  _T_76 = 5'h6 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_77 = _T_76 ? {{1'd0}, _T_49} : _T_75; // @[Mux.scala 68:16]
  wire  _T_78 = 5'h5 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_79 = _T_78 ? {{1'd0}, _T_45} : _T_77; // @[Mux.scala 68:16]
  wire  _T_80 = 5'h4 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_81 = _T_80 ? {{1'd0}, _T_41} : _T_79; // @[Mux.scala 68:16]
  wire  _T_82 = 5'h3 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_83 = _T_82 ? {{1'd0}, _T_37} : _T_81; // @[Mux.scala 68:16]
  wire  _T_84 = 5'h2 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_85 = _T_84 ? {{1'd0}, _T_33} : _T_83; // @[Mux.scala 68:16]
  wire  _T_86 = 5'h1 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] _T_87 = _T_86 ? {{1'd0}, _T_29} : _T_85; // @[Mux.scala 68:16]
  wire  _T_88 = 5'h0 == io_fu_in_bits_ops_fu_op; // @[Mux.scala 68:19]
  wire [34:0] br_info = _T_88 ? {{1'd0}, _T_26} : _T_87; // @[Mux.scala 68:16]
  assign io_fu_out_valid = io_fu_in_valid & br_info[33]; // @[bru.scala 42:19]
  assign io_fu_out_bits_wb_v = br_info[32]; // @[bru.scala 43:21 bru.scala 44:23]
  assign io_fu_out_bits_wb_pc = io_fu_in_bits_wb_pc; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[bru.scala 43:21]
  assign io_fu_out_bits_wb_wen = br_info[32]; // @[bru.scala 43:21 bru.scala 45:25]
  assign io_fu_out_bits_wb_data = io_fu_in_bits_wb_pc + 32'h8; // @[bru.scala 43:21 bru.scala 46:26]
  assign io_fu_out_bits_wb_is_ds = io_fu_in_bits_wb_is_ds; // @[bru.scala 43:21]
  assign io_fu_out_bits_br_target = br_info[31:0]; // @[bru.scala 48:28]
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input  [31:0] io_fu_in_bits_pc,
  input  [5:0]  io_fu_in_bits_instr_op,
  input  [4:0]  io_fu_in_bits_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_instr_shamt,
  input  [5:0]  io_fu_in_bits_instr_func,
  input  [2:0]  io_fu_in_bits_fu_type,
  input  [4:0]  io_fu_in_bits_fu_op,
  input  [1:0]  io_fu_in_bits_op1_sel,
  input  [2:0]  io_fu_in_bits_op2_sel,
  input  [1:0]  io_fu_in_bits_opd_sel,
  input  [4:0]  io_fu_in_bits_ex_et,
  input  [4:0]  io_fu_in_bits_ex_code,
  input  [31:0] io_fu_in_bits_ex_addr,
  input  [7:0]  io_fu_in_bits_ex_asid,
  input         io_fu_out_ready,
  output        io_fu_out_valid,
  output        io_fu_out_bits_wb_v,
  output [7:0]  io_fu_out_bits_wb_id,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output [4:0]  io_fu_out_bits_wb_rd_idx,
  output        io_fu_out_bits_wb_wen,
  output [31:0] io_fu_out_bits_wb_data,
  output        io_fu_out_bits_wb_is_ds,
  output        io_fu_out_bits_wb_is_br,
  output [31:0] io_fu_out_bits_wb_npc,
  output [2:0]  io_fu_out_bits_ops_fu_type,
  output [4:0]  io_fu_out_bits_ops_fu_op,
  output [31:0] io_fu_out_bits_ops_op1,
  output [31:0] io_fu_out_bits_ops_op2,
  output [4:0]  io_fu_out_bits_ex_et,
  output [4:0]  io_fu_out_bits_ex_code,
  output [31:0] io_fu_out_bits_ex_addr,
  output [7:0]  io_fu_out_bits_ex_asid,
  output        io_br_flush_valid,
  output [31:0] io_br_flush_bits_br_target,
  output [4:0]  io_rfio_rs_idx,
  output [4:0]  io_rfio_rt_idx,
  output        io_rfio_wen,
  output [7:0]  io_rfio_wid,
  output [4:0]  io_rfio_rd_idx,
  input         io_rfio_rs_data_valid,
  input  [31:0] io_rfio_rs_data_bits,
  input         io_rfio_rt_data_valid,
  input  [31:0] io_rfio_rt_data_bits
);
  wire  bru_io_fu_in_valid; // @[isu.scala 22:19]
  wire [31:0] bru_io_fu_in_bits_wb_pc; // @[isu.scala 22:19]
  wire [5:0] bru_io_fu_in_bits_wb_instr_op; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_in_bits_wb_instr_rs_idx; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_in_bits_wb_instr_rt_idx; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_in_bits_wb_instr_rd_idx; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_in_bits_wb_instr_shamt; // @[isu.scala 22:19]
  wire [5:0] bru_io_fu_in_bits_wb_instr_func; // @[isu.scala 22:19]
  wire  bru_io_fu_in_bits_wb_is_ds; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_in_bits_ops_fu_op; // @[isu.scala 22:19]
  wire [31:0] bru_io_fu_in_bits_ops_op1; // @[isu.scala 22:19]
  wire [31:0] bru_io_fu_in_bits_ops_op2; // @[isu.scala 22:19]
  wire  bru_io_fu_out_valid; // @[isu.scala 22:19]
  wire  bru_io_fu_out_bits_wb_v; // @[isu.scala 22:19]
  wire [31:0] bru_io_fu_out_bits_wb_pc; // @[isu.scala 22:19]
  wire [5:0] bru_io_fu_out_bits_wb_instr_op; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_out_bits_wb_instr_rs_idx; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_out_bits_wb_instr_rt_idx; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_out_bits_wb_instr_rd_idx; // @[isu.scala 22:19]
  wire [4:0] bru_io_fu_out_bits_wb_instr_shamt; // @[isu.scala 22:19]
  wire [5:0] bru_io_fu_out_bits_wb_instr_func; // @[isu.scala 22:19]
  wire  bru_io_fu_out_bits_wb_wen; // @[isu.scala 22:19]
  wire [31:0] bru_io_fu_out_bits_wb_data; // @[isu.scala 22:19]
  wire  bru_io_fu_out_bits_wb_is_ds; // @[isu.scala 22:19]
  wire [31:0] bru_io_fu_out_bits_br_target; // @[isu.scala 22:19]
  reg [7:0] instr_id; // @[isu.scala 26:25]
  reg [31:0] _RAND_0;
  wire  _T = io_fu_out_ready & io_fu_out_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_2 = instr_id + 8'h1; // @[isu.scala 27:50]
  wire  _T_4 = io_fu_in_bits_opd_sel != 2'h0; // @[isu.scala 32:60]
  wire  _T_6 = 2'h3 == io_fu_in_bits_opd_sel; // @[Mux.scala 68:19]
  wire [4:0] _T_7 = _T_6 ? 5'h1f : 5'h0; // @[Mux.scala 68:16]
  wire  _T_8 = 2'h2 == io_fu_in_bits_opd_sel; // @[Mux.scala 68:19]
  wire [4:0] _T_9 = _T_8 ? io_fu_in_bits_instr_rt_idx : _T_7; // @[Mux.scala 68:16]
  wire  _T_10 = 2'h1 == io_fu_in_bits_opd_sel; // @[Mux.scala 68:19]
  wire  _T_12 = io_fu_in_bits_op1_sel == 2'h1; // @[isu.scala 40:45]
  wire  _T_13 = io_fu_in_bits_op1_sel == 2'h3; // @[isu.scala 41:28]
  wire  _T_14 = _T_12 | _T_13; // @[isu.scala 40:57]
  wire  _T_15 = io_fu_in_bits_op2_sel == 3'h1; // @[isu.scala 42:28]
  wire  _T_16 = _T_14 | _T_15; // @[isu.scala 41:41]
  wire  rs_ready = _T_16 ? io_rfio_rs_data_valid : 1'h1; // @[isu.scala 40:21]
  wire  _T_17 = io_fu_in_bits_op1_sel == 2'h2; // @[isu.scala 44:45]
  wire  _T_18 = io_fu_in_bits_op2_sel == 3'h2; // @[isu.scala 45:28]
  wire  _T_19 = _T_17 | _T_18; // @[isu.scala 44:57]
  wire  rt_ready = _T_19 ? io_rfio_rt_data_valid : 1'h1; // @[isu.scala 44:21]
  wire  reg_ready = rs_ready & rt_ready; // @[isu.scala 47:28]
  wire [15:0] _T_21 = {io_fu_in_bits_instr_rd_idx,io_fu_in_bits_instr_shamt,io_fu_in_bits_instr_func}; // @[Cat.scala 29:58]
  wire [15:0] _T_23 = {io_fu_in_bits_instr_rd_idx,io_fu_in_bits_instr_shamt,io_fu_in_bits_instr_func}; // @[isu.scala 51:34]
  wire [31:0] se_imm = {{16{_T_23[15]}},_T_23}; // @[isu.scala 51:56]
  wire [31:0] ue_imm = {io_fu_in_bits_instr_rd_idx,io_fu_in_bits_instr_shamt,io_fu_in_bits_instr_func,16'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_34 = io_rfio_rs_data_bits + se_imm; // @[isu.scala 60:53]
  wire [31:0] _T_35 = _T_12 ? io_rfio_rs_data_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_36 = _T_17 ? io_rfio_rt_data_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_37 = _T_13 ? _T_34 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_38 = _T_35 | _T_36; // @[Mux.scala 27:72]
  wire  _T_42 = io_fu_in_bits_op2_sel == 3'h3; // @[isu.scala 66:28]
  wire  _T_43 = io_fu_in_bits_op2_sel == 3'h4; // @[isu.scala 67:28]
  wire  _T_44 = io_fu_in_bits_op2_sel == 3'h5; // @[isu.scala 68:28]
  wire  _T_45 = io_fu_in_bits_op2_sel == 3'h6; // @[isu.scala 69:28]
  wire  _T_46 = io_fu_in_bits_op2_sel == 3'h7; // @[isu.scala 70:28]
  wire [31:0] _T_47 = _T_15 ? io_rfio_rs_data_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_48 = _T_18 ? io_rfio_rt_data_bits : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_49 = _T_42 ? se_imm : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_50 = _T_43 ? ue_imm : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] ze_imm = {{16'd0}, _T_21}; // @[isu.scala 52:34 isu.scala 52:34]
  wire [31:0] _T_51 = _T_44 ? ze_imm : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] shamt_ext = {{27'd0}, io_fu_in_bits_instr_shamt}; // @[isu.scala 50:39 isu.scala 50:39]
  wire [31:0] _T_52 = _T_45 ? shamt_ext : 32'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_53 = _T_46 ? io_fu_in_bits_instr_rt_idx : 5'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_54 = _T_47 | _T_48; // @[Mux.scala 27:72]
  wire [31:0] _T_55 = _T_54 | _T_49; // @[Mux.scala 27:72]
  wire [31:0] _T_56 = _T_55 | _T_50; // @[Mux.scala 27:72]
  wire [31:0] _T_57 = _T_56 | _T_51; // @[Mux.scala 27:72]
  wire [31:0] _T_58 = _T_57 | _T_52; // @[Mux.scala 27:72]
  wire [31:0] _GEN_4 = {{27'd0}, _T_53}; // @[Mux.scala 27:72]
  reg  is_delayslot; // @[isu.scala 73:29]
  reg [31:0] _RAND_1;
  reg [31:0] br_target; // @[isu.scala 74:26]
  reg [31:0] _RAND_2;
  wire  _T_62 = io_fu_in_bits_fu_type == 3'h2; // @[isu.scala 76:51]
  wire  _T_63 = _T & _T_62; // @[isu.scala 76:26]
  wire [31:0] _T_65 = io_fu_out_bits_wb_pc + 32'h8; // @[isu.scala 80:28]
  wire  _GEN_1 = _T ? 1'h0 : is_delayslot; // @[isu.scala 81:34]
  wire  _GEN_2 = _T_63 | _GEN_1; // @[isu.scala 76:63]
  wire [31:0] _T_74 = io_fu_out_bits_wb_pc + 32'h4; // @[isu.scala 96:26]
  BRU bru ( // @[isu.scala 22:19]
    .io_fu_in_valid(bru_io_fu_in_valid),
    .io_fu_in_bits_wb_pc(bru_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(bru_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(bru_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(bru_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(bru_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(bru_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(bru_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_is_ds(bru_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_ops_fu_op(bru_io_fu_in_bits_ops_fu_op),
    .io_fu_in_bits_ops_op1(bru_io_fu_in_bits_ops_op1),
    .io_fu_in_bits_ops_op2(bru_io_fu_in_bits_ops_op2),
    .io_fu_out_valid(bru_io_fu_out_valid),
    .io_fu_out_bits_wb_v(bru_io_fu_out_bits_wb_v),
    .io_fu_out_bits_wb_pc(bru_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(bru_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(bru_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(bru_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(bru_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(bru_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(bru_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_wen(bru_io_fu_out_bits_wb_wen),
    .io_fu_out_bits_wb_data(bru_io_fu_out_bits_wb_data),
    .io_fu_out_bits_wb_is_ds(bru_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_br_target(bru_io_fu_out_bits_br_target)
  );
  assign io_fu_in_ready = io_fu_out_ready & reg_ready; // @[isu.scala 87:18]
  assign io_fu_out_valid = io_fu_in_valid & reg_ready; // @[isu.scala 88:19]
  assign io_fu_out_bits_wb_v = _T_62 & bru_io_fu_out_bits_wb_v; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_id = instr_id; // @[isu.scala 93:21 isu.scala 97:24]
  assign io_fu_out_bits_wb_pc = _T_62 ? bru_io_fu_out_bits_wb_pc : io_fu_in_bits_pc; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_instr_op = _T_62 ? bru_io_fu_out_bits_wb_instr_op : io_fu_in_bits_instr_op; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_instr_rs_idx = _T_62 ? bru_io_fu_out_bits_wb_instr_rs_idx : io_fu_in_bits_instr_rs_idx; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_instr_rt_idx = _T_62 ? bru_io_fu_out_bits_wb_instr_rt_idx : io_fu_in_bits_instr_rt_idx; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_instr_rd_idx = _T_62 ? bru_io_fu_out_bits_wb_instr_rd_idx : io_fu_in_bits_instr_rd_idx; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_instr_shamt = _T_62 ? bru_io_fu_out_bits_wb_instr_shamt : io_fu_in_bits_instr_shamt; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_instr_func = _T_62 ? bru_io_fu_out_bits_wb_instr_func : io_fu_in_bits_instr_func; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_rd_idx = io_rfio_rd_idx; // @[isu.scala 93:21 isu.scala 98:28]
  assign io_fu_out_bits_wb_wen = _T_62 & bru_io_fu_out_bits_wb_wen; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_data = _T_62 ? bru_io_fu_out_bits_wb_data : 32'h0; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_is_ds = _T_62 ? bru_io_fu_out_bits_wb_is_ds : is_delayslot; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_is_br = io_fu_in_bits_fu_type == 3'h2; // @[isu.scala 93:21]
  assign io_fu_out_bits_wb_npc = is_delayslot ? br_target : _T_74; // @[isu.scala 93:21 isu.scala 95:25]
  assign io_fu_out_bits_ops_fu_type = io_fu_in_bits_fu_type; // @[isu.scala 89:30]
  assign io_fu_out_bits_ops_fu_op = io_fu_in_bits_fu_op; // @[isu.scala 90:28]
  assign io_fu_out_bits_ops_op1 = _T_38 | _T_37; // @[isu.scala 91:26]
  assign io_fu_out_bits_ops_op2 = _T_58 | _GEN_4; // @[isu.scala 92:26]
  assign io_fu_out_bits_ex_et = io_fu_in_bits_ex_et; // @[isu.scala 99:21]
  assign io_fu_out_bits_ex_code = io_fu_in_bits_ex_code; // @[isu.scala 99:21]
  assign io_fu_out_bits_ex_addr = io_fu_in_bits_ex_addr; // @[isu.scala 99:21]
  assign io_fu_out_bits_ex_asid = io_fu_in_bits_ex_asid; // @[isu.scala 99:21]
  assign io_br_flush_valid = bru_io_fu_out_valid & _T; // @[isu.scala 106:21]
  assign io_br_flush_bits_br_target = bru_io_fu_out_bits_br_target; // @[isu.scala 107:30]
  assign io_rfio_rs_idx = io_fu_in_bits_instr_rs_idx; // @[isu.scala 30:18]
  assign io_rfio_rt_idx = io_fu_in_bits_instr_rt_idx; // @[isu.scala 31:18]
  assign io_rfio_wen = _T & _T_4; // @[isu.scala 32:15]
  assign io_rfio_wid = instr_id; // @[isu.scala 33:15]
  assign io_rfio_rd_idx = _T_10 ? io_fu_in_bits_instr_rd_idx : _T_9; // @[isu.scala 34:18]
  assign bru_io_fu_in_valid = io_fu_in_valid & _T_62; // @[isu.scala 102:22]
  assign bru_io_fu_in_bits_wb_pc = io_fu_in_bits_pc; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_instr_op = io_fu_in_bits_instr_op; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_instr_rs_idx = io_fu_in_bits_instr_rs_idx; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_instr_rt_idx = io_fu_in_bits_instr_rt_idx; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_instr_rd_idx = io_fu_in_bits_instr_rd_idx; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_instr_shamt = io_fu_in_bits_instr_shamt; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_instr_func = io_fu_in_bits_instr_func; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_wb_is_ds = is_delayslot; // @[isu.scala 103:24]
  assign bru_io_fu_in_bits_ops_fu_op = io_fu_out_bits_ops_fu_op; // @[isu.scala 104:25]
  assign bru_io_fu_in_bits_ops_op1 = io_fu_out_bits_ops_op1; // @[isu.scala 104:25]
  assign bru_io_fu_in_bits_ops_op2 = io_fu_out_bits_ops_op2; // @[isu.scala 104:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  instr_id = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  is_delayslot = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  br_target = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      instr_id <= 8'h0;
    end else if (_T) begin
      instr_id <= _T_2;
    end
    if (reset) begin
      is_delayslot <= 1'h0;
    end else begin
      is_delayslot <= _GEN_2;
    end
    if (reset) begin
      br_target <= 32'h0;
    end else if (_T_63) begin
      if (io_br_flush_valid) begin
        br_target <= io_br_flush_bits_br_target;
      end else begin
        br_target <= _T_65;
      end
    end
  end
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input  [31:0] io_fu_in_bits_pc,
  input  [31:0] io_fu_in_bits_instr,
  input  [4:0]  io_fu_in_bits_ex_et,
  input  [4:0]  io_fu_in_bits_ex_code,
  input  [31:0] io_fu_in_bits_ex_addr,
  input  [7:0]  io_fu_in_bits_ex_asid,
  input         io_fu_out_ready,
  output        io_fu_out_valid,
  output        io_fu_out_bits_wb_v,
  output [7:0]  io_fu_out_bits_wb_id,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output [4:0]  io_fu_out_bits_wb_rd_idx,
  output        io_fu_out_bits_wb_wen,
  output [31:0] io_fu_out_bits_wb_data,
  output        io_fu_out_bits_wb_is_ds,
  output        io_fu_out_bits_wb_is_br,
  output [31:0] io_fu_out_bits_wb_npc,
  output [2:0]  io_fu_out_bits_ops_fu_type,
  output [4:0]  io_fu_out_bits_ops_fu_op,
  output [31:0] io_fu_out_bits_ops_op1,
  output [31:0] io_fu_out_bits_ops_op2,
  output [4:0]  io_fu_out_bits_ex_et,
  output [4:0]  io_fu_out_bits_ex_code,
  output [31:0] io_fu_out_bits_ex_addr,
  output [7:0]  io_fu_out_bits_ex_asid,
  output        io_br_flush_valid,
  output [31:0] io_br_flush_bits_br_target,
  output [4:0]  io_rfio_rs_idx,
  output [4:0]  io_rfio_rt_idx,
  output        io_rfio_wen,
  output [7:0]  io_rfio_wid,
  output [4:0]  io_rfio_rd_idx,
  input         io_rfio_rs_data_valid,
  input  [31:0] io_rfio_rs_data_bits,
  input         io_rfio_rt_data_valid,
  input  [31:0] io_rfio_rt_data_bits,
  input         io_ex_flush_valid
);
  wire  isu_clock; // @[idu.scala 21:19]
  wire  isu_reset; // @[idu.scala 21:19]
  wire  isu_io_fu_in_ready; // @[idu.scala 21:19]
  wire  isu_io_fu_in_valid; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_in_bits_pc; // @[idu.scala 21:19]
  wire [5:0] isu_io_fu_in_bits_instr_op; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_instr_rs_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_instr_rt_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_instr_rd_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_instr_shamt; // @[idu.scala 21:19]
  wire [5:0] isu_io_fu_in_bits_instr_func; // @[idu.scala 21:19]
  wire [2:0] isu_io_fu_in_bits_fu_type; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_fu_op; // @[idu.scala 21:19]
  wire [1:0] isu_io_fu_in_bits_op1_sel; // @[idu.scala 21:19]
  wire [2:0] isu_io_fu_in_bits_op2_sel; // @[idu.scala 21:19]
  wire [1:0] isu_io_fu_in_bits_opd_sel; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_ex_et; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_in_bits_ex_code; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_in_bits_ex_addr; // @[idu.scala 21:19]
  wire [7:0] isu_io_fu_in_bits_ex_asid; // @[idu.scala 21:19]
  wire  isu_io_fu_out_ready; // @[idu.scala 21:19]
  wire  isu_io_fu_out_valid; // @[idu.scala 21:19]
  wire  isu_io_fu_out_bits_wb_v; // @[idu.scala 21:19]
  wire [7:0] isu_io_fu_out_bits_wb_id; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_out_bits_wb_pc; // @[idu.scala 21:19]
  wire [5:0] isu_io_fu_out_bits_wb_instr_op; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_wb_instr_rs_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_wb_instr_rt_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_wb_instr_rd_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_wb_instr_shamt; // @[idu.scala 21:19]
  wire [5:0] isu_io_fu_out_bits_wb_instr_func; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_wb_rd_idx; // @[idu.scala 21:19]
  wire  isu_io_fu_out_bits_wb_wen; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_out_bits_wb_data; // @[idu.scala 21:19]
  wire  isu_io_fu_out_bits_wb_is_ds; // @[idu.scala 21:19]
  wire  isu_io_fu_out_bits_wb_is_br; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_out_bits_wb_npc; // @[idu.scala 21:19]
  wire [2:0] isu_io_fu_out_bits_ops_fu_type; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_ops_fu_op; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_out_bits_ops_op1; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_out_bits_ops_op2; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_ex_et; // @[idu.scala 21:19]
  wire [4:0] isu_io_fu_out_bits_ex_code; // @[idu.scala 21:19]
  wire [31:0] isu_io_fu_out_bits_ex_addr; // @[idu.scala 21:19]
  wire [7:0] isu_io_fu_out_bits_ex_asid; // @[idu.scala 21:19]
  wire  isu_io_br_flush_valid; // @[idu.scala 21:19]
  wire [31:0] isu_io_br_flush_bits_br_target; // @[idu.scala 21:19]
  wire [4:0] isu_io_rfio_rs_idx; // @[idu.scala 21:19]
  wire [4:0] isu_io_rfio_rt_idx; // @[idu.scala 21:19]
  wire  isu_io_rfio_wen; // @[idu.scala 21:19]
  wire [7:0] isu_io_rfio_wid; // @[idu.scala 21:19]
  wire [4:0] isu_io_rfio_rd_idx; // @[idu.scala 21:19]
  wire  isu_io_rfio_rs_data_valid; // @[idu.scala 21:19]
  wire [31:0] isu_io_rfio_rs_data_bits; // @[idu.scala 21:19]
  wire  isu_io_rfio_rt_data_valid; // @[idu.scala 21:19]
  wire [31:0] isu_io_rfio_rt_data_bits; // @[idu.scala 21:19]
  wire  _T_30 = io_fu_in_ready & io_fu_in_valid; // @[Decoupled.scala 40:37]
  reg [31:0] fu_in_pc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_0;
  reg [31:0] fu_in_instr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [4:0] fu_in_ex_et; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [4:0] fu_in_ex_code; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [31:0] fu_in_ex_addr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [7:0] fu_in_ex_asid; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg  fu_valid; // @[idu.scala 23:25]
  reg [31:0] _RAND_6;
  wire  _T_32 = ~fu_valid; // @[idu.scala 26:21]
  wire [31:0] _T_34 = fu_in_instr & 32'hffe00000; // @[Lookup.scala 31:38]
  wire  _T_35 = 32'h3c000000 == _T_34; // @[Lookup.scala 31:38]
  wire [31:0] _T_36 = fu_in_instr & 32'hfc0007ff; // @[Lookup.scala 31:38]
  wire  _T_37 = 32'h20 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_39 = 32'h21 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_41 = 32'h22 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_43 = 32'h23 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_45 = 32'h2a == _T_36; // @[Lookup.scala 31:38]
  wire  _T_47 = 32'h2b == _T_36; // @[Lookup.scala 31:38]
  wire  _T_49 = 32'h24 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_51 = 32'h25 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_53 = 32'h26 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_55 = 32'h27 == _T_36; // @[Lookup.scala 31:38]
  wire [31:0] _T_56 = fu_in_instr & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _T_57 = 32'h28000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_59 = 32'h2c000000 == _T_56; // @[Lookup.scala 31:38]
  wire [31:0] _T_60 = fu_in_instr & 32'hffe0003f; // @[Lookup.scala 31:38]
  wire  _T_61 = 32'h0 == _T_60; // @[Lookup.scala 31:38]
  wire  _T_63 = 32'h3 == _T_60; // @[Lookup.scala 31:38]
  wire  _T_65 = 32'h2 == _T_60; // @[Lookup.scala 31:38]
  wire  _T_67 = 32'h7 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_69 = 32'h6 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_71 = 32'h4 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_73 = 32'h20000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_75 = 32'h24000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_77 = 32'h30000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_79 = 32'h34000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_81 = 32'h38000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_83 = 32'hb == _T_36; // @[Lookup.scala 31:38]
  wire  _T_85 = 32'ha == _T_36; // @[Lookup.scala 31:38]
  wire  _T_87 = 32'h70000020 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_89 = 32'h70000021 == _T_36; // @[Lookup.scala 31:38]
  wire [31:0] _T_90 = fu_in_instr & 32'hffe007ff; // @[Lookup.scala 31:38]
  wire  _T_91 = 32'h7c000420 == _T_90; // @[Lookup.scala 31:38]
  wire  _T_93 = 32'h7c000620 == _T_90; // @[Lookup.scala 31:38]
  wire  _T_95 = 32'h7c0000a0 == _T_36; // @[Lookup.scala 31:38]
  wire [31:0] _T_96 = fu_in_instr & 32'hfc00003f; // @[Lookup.scala 31:38]
  wire  _T_97 = 32'h7c000004 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_99 = 32'h7c000000 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_101 = 32'h200002 == _T_60; // @[Lookup.scala 31:38]
  wire  _T_103 = 32'h46 == _T_36; // @[Lookup.scala 31:38]
  wire  _T_105 = 32'h10000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_107 = 32'h14000000 == _T_56; // @[Lookup.scala 31:38]
  wire [31:0] _T_108 = fu_in_instr & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _T_109 = 32'h18000000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_111 = 32'h4010000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_113 = 32'h4000000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_115 = 32'h1c000000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_117 = 32'h4110000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_119 = 32'h4100000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_121 = 32'h8000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_123 = 32'hc000000 == _T_56; // @[Lookup.scala 31:38]
  wire [31:0] _T_124 = fu_in_instr & 32'hfc1ff83f; // @[Lookup.scala 31:38]
  wire  _T_125 = 32'h8 == _T_124; // @[Lookup.scala 31:38]
  wire  _T_127 = 32'h9 == _T_36; // @[Lookup.scala 31:38]
  wire [31:0] _T_128 = fu_in_instr & 32'hffff07ff; // @[Lookup.scala 31:38]
  wire  _T_129 = 32'h10 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 32'h12 == _T_128; // @[Lookup.scala 31:38]
  wire [31:0] _T_132 = fu_in_instr & 32'hfc1fffff; // @[Lookup.scala 31:38]
  wire  _T_133 = 32'h11 == _T_132; // @[Lookup.scala 31:38]
  wire  _T_135 = 32'h13 == _T_132; // @[Lookup.scala 31:38]
  wire  _T_137 = 32'h70000002 == _T_36; // @[Lookup.scala 31:38]
  wire [31:0] _T_138 = fu_in_instr & 32'hfc00ffff; // @[Lookup.scala 31:38]
  wire  _T_139 = 32'h18 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_141 = 32'h19 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_143 = 32'h1a == _T_138; // @[Lookup.scala 31:38]
  wire  _T_145 = 32'h1b == _T_138; // @[Lookup.scala 31:38]
  wire  _T_147 = 32'h70000000 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_149 = 32'h70000001 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_151 = 32'h70000004 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_153 = 32'h70000005 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_155 = 32'h8c000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_157 = 32'h84000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_159 = 32'h94000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_161 = 32'h80000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_163 = 32'h90000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_165 = 32'h88000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_167 = 32'h98000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_169 = 32'hac000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_171 = 32'ha4000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_173 = 32'ha0000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_175 = 32'ha8000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_177 = 32'hb8000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_179 = 32'hc0000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_181 = 32'he0000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_183 = 32'hc == _T_96; // @[Lookup.scala 31:38]
  wire  _T_185 = 32'hd == _T_96; // @[Lookup.scala 31:38]
  wire  _T_187 = 32'h42000018 == fu_in_instr; // @[Lookup.scala 31:38]
  wire [31:0] _T_188 = fu_in_instr & 32'hffe007f8; // @[Lookup.scala 31:38]
  wire  _T_189 = 32'h40000000 == _T_188; // @[Lookup.scala 31:38]
  wire  _T_191 = 32'h40800000 == _T_188; // @[Lookup.scala 31:38]
  wire  _T_193 = 32'hbc000000 == _T_56; // @[Lookup.scala 31:38]
  wire [31:0] _T_194 = fu_in_instr & 32'hfffff83f; // @[Lookup.scala 31:38]
  wire  _T_195 = 32'hf == _T_194; // @[Lookup.scala 31:38]
  wire  _T_197 = 32'hcc000000 == _T_56; // @[Lookup.scala 31:38]
  wire  _T_199 = 32'h42000008 == fu_in_instr; // @[Lookup.scala 31:38]
  wire  _T_201 = 32'h42000001 == fu_in_instr; // @[Lookup.scala 31:38]
  wire  _T_203 = 32'h42000002 == fu_in_instr; // @[Lookup.scala 31:38]
  wire  _T_205 = 32'h42000006 == fu_in_instr; // @[Lookup.scala 31:38]
  wire  _T_207 = 32'h30 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_209 = 32'h31 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_211 = 32'h32 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_213 = 32'h33 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_215 = 32'h34 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_217 = 32'h36 == _T_96; // @[Lookup.scala 31:38]
  wire  _T_219 = 32'h4080000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_221 = 32'h4090000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_223 = 32'h40a0000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_225 = 32'h40b0000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_227 = 32'h40c0000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_229 = 32'h40e0000 == _T_108; // @[Lookup.scala 31:38]
  wire  _T_231 = _T_227 | _T_229; // @[Lookup.scala 33:37]
  wire  _T_232 = _T_225 | _T_231; // @[Lookup.scala 33:37]
  wire  _T_233 = _T_223 | _T_232; // @[Lookup.scala 33:37]
  wire  _T_234 = _T_221 | _T_233; // @[Lookup.scala 33:37]
  wire  _T_235 = _T_219 | _T_234; // @[Lookup.scala 33:37]
  wire  _T_236 = _T_217 | _T_235; // @[Lookup.scala 33:37]
  wire  _T_237 = _T_215 | _T_236; // @[Lookup.scala 33:37]
  wire  _T_238 = _T_213 | _T_237; // @[Lookup.scala 33:37]
  wire  _T_239 = _T_211 | _T_238; // @[Lookup.scala 33:37]
  wire  _T_240 = _T_209 | _T_239; // @[Lookup.scala 33:37]
  wire  _T_241 = _T_207 | _T_240; // @[Lookup.scala 33:37]
  wire  _T_242 = _T_205 | _T_241; // @[Lookup.scala 33:37]
  wire  _T_243 = _T_203 | _T_242; // @[Lookup.scala 33:37]
  wire  _T_244 = _T_201 | _T_243; // @[Lookup.scala 33:37]
  wire  _T_245 = _T_199 | _T_244; // @[Lookup.scala 33:37]
  wire  _T_246 = _T_197 | _T_245; // @[Lookup.scala 33:37]
  wire  _T_247 = _T_195 | _T_246; // @[Lookup.scala 33:37]
  wire  _T_248 = _T_193 | _T_247; // @[Lookup.scala 33:37]
  wire  _T_249 = _T_191 | _T_248; // @[Lookup.scala 33:37]
  wire  _T_250 = _T_189 | _T_249; // @[Lookup.scala 33:37]
  wire  _T_251 = _T_187 | _T_250; // @[Lookup.scala 33:37]
  wire  _T_252 = _T_185 | _T_251; // @[Lookup.scala 33:37]
  wire  _T_253 = _T_183 | _T_252; // @[Lookup.scala 33:37]
  wire  _T_254 = _T_181 | _T_253; // @[Lookup.scala 33:37]
  wire  _T_255 = _T_179 | _T_254; // @[Lookup.scala 33:37]
  wire  _T_256 = _T_177 | _T_255; // @[Lookup.scala 33:37]
  wire  _T_257 = _T_175 | _T_256; // @[Lookup.scala 33:37]
  wire  _T_258 = _T_173 | _T_257; // @[Lookup.scala 33:37]
  wire  _T_259 = _T_171 | _T_258; // @[Lookup.scala 33:37]
  wire  _T_260 = _T_169 | _T_259; // @[Lookup.scala 33:37]
  wire  _T_261 = _T_167 | _T_260; // @[Lookup.scala 33:37]
  wire  _T_262 = _T_165 | _T_261; // @[Lookup.scala 33:37]
  wire  _T_263 = _T_163 | _T_262; // @[Lookup.scala 33:37]
  wire  _T_264 = _T_161 | _T_263; // @[Lookup.scala 33:37]
  wire  _T_265 = _T_159 | _T_264; // @[Lookup.scala 33:37]
  wire  _T_266 = _T_157 | _T_265; // @[Lookup.scala 33:37]
  wire  _T_267 = _T_155 | _T_266; // @[Lookup.scala 33:37]
  wire  _T_268 = _T_153 | _T_267; // @[Lookup.scala 33:37]
  wire  _T_269 = _T_151 | _T_268; // @[Lookup.scala 33:37]
  wire  _T_270 = _T_149 | _T_269; // @[Lookup.scala 33:37]
  wire  _T_271 = _T_147 | _T_270; // @[Lookup.scala 33:37]
  wire  _T_272 = _T_145 | _T_271; // @[Lookup.scala 33:37]
  wire  _T_273 = _T_143 | _T_272; // @[Lookup.scala 33:37]
  wire  _T_274 = _T_141 | _T_273; // @[Lookup.scala 33:37]
  wire  _T_275 = _T_139 | _T_274; // @[Lookup.scala 33:37]
  wire  _T_276 = _T_137 | _T_275; // @[Lookup.scala 33:37]
  wire  _T_277 = _T_135 | _T_276; // @[Lookup.scala 33:37]
  wire  _T_278 = _T_133 | _T_277; // @[Lookup.scala 33:37]
  wire  _T_279 = _T_131 | _T_278; // @[Lookup.scala 33:37]
  wire  _T_280 = _T_129 | _T_279; // @[Lookup.scala 33:37]
  wire  _T_281 = _T_127 | _T_280; // @[Lookup.scala 33:37]
  wire  _T_282 = _T_125 | _T_281; // @[Lookup.scala 33:37]
  wire  _T_283 = _T_123 | _T_282; // @[Lookup.scala 33:37]
  wire  _T_284 = _T_121 | _T_283; // @[Lookup.scala 33:37]
  wire  _T_285 = _T_119 | _T_284; // @[Lookup.scala 33:37]
  wire  _T_286 = _T_117 | _T_285; // @[Lookup.scala 33:37]
  wire  _T_287 = _T_115 | _T_286; // @[Lookup.scala 33:37]
  wire  _T_288 = _T_113 | _T_287; // @[Lookup.scala 33:37]
  wire  _T_289 = _T_111 | _T_288; // @[Lookup.scala 33:37]
  wire  _T_290 = _T_109 | _T_289; // @[Lookup.scala 33:37]
  wire  _T_291 = _T_107 | _T_290; // @[Lookup.scala 33:37]
  wire  _T_292 = _T_105 | _T_291; // @[Lookup.scala 33:37]
  wire  _T_293 = _T_103 | _T_292; // @[Lookup.scala 33:37]
  wire  _T_294 = _T_101 | _T_293; // @[Lookup.scala 33:37]
  wire  _T_295 = _T_99 | _T_294; // @[Lookup.scala 33:37]
  wire  _T_296 = _T_97 | _T_295; // @[Lookup.scala 33:37]
  wire  _T_297 = _T_95 | _T_296; // @[Lookup.scala 33:37]
  wire  _T_298 = _T_93 | _T_297; // @[Lookup.scala 33:37]
  wire  _T_299 = _T_91 | _T_298; // @[Lookup.scala 33:37]
  wire  _T_300 = _T_89 | _T_299; // @[Lookup.scala 33:37]
  wire  _T_301 = _T_87 | _T_300; // @[Lookup.scala 33:37]
  wire  _T_302 = _T_85 | _T_301; // @[Lookup.scala 33:37]
  wire  _T_303 = _T_83 | _T_302; // @[Lookup.scala 33:37]
  wire  _T_304 = _T_81 | _T_303; // @[Lookup.scala 33:37]
  wire  _T_305 = _T_79 | _T_304; // @[Lookup.scala 33:37]
  wire  _T_306 = _T_77 | _T_305; // @[Lookup.scala 33:37]
  wire  _T_307 = _T_75 | _T_306; // @[Lookup.scala 33:37]
  wire  _T_308 = _T_73 | _T_307; // @[Lookup.scala 33:37]
  wire  _T_309 = _T_71 | _T_308; // @[Lookup.scala 33:37]
  wire  _T_310 = _T_69 | _T_309; // @[Lookup.scala 33:37]
  wire  _T_311 = _T_67 | _T_310; // @[Lookup.scala 33:37]
  wire  _T_312 = _T_65 | _T_311; // @[Lookup.scala 33:37]
  wire  _T_313 = _T_63 | _T_312; // @[Lookup.scala 33:37]
  wire  _T_314 = _T_61 | _T_313; // @[Lookup.scala 33:37]
  wire  _T_315 = _T_59 | _T_314; // @[Lookup.scala 33:37]
  wire  _T_316 = _T_57 | _T_315; // @[Lookup.scala 33:37]
  wire  _T_317 = _T_55 | _T_316; // @[Lookup.scala 33:37]
  wire  _T_318 = _T_53 | _T_317; // @[Lookup.scala 33:37]
  wire  _T_319 = _T_51 | _T_318; // @[Lookup.scala 33:37]
  wire  _T_320 = _T_49 | _T_319; // @[Lookup.scala 33:37]
  wire  _T_321 = _T_47 | _T_320; // @[Lookup.scala 33:37]
  wire  _T_322 = _T_45 | _T_321; // @[Lookup.scala 33:37]
  wire  _T_323 = _T_43 | _T_322; // @[Lookup.scala 33:37]
  wire  _T_324 = _T_41 | _T_323; // @[Lookup.scala 33:37]
  wire  _T_325 = _T_39 | _T_324; // @[Lookup.scala 33:37]
  wire  _T_326 = _T_37 | _T_325; // @[Lookup.scala 33:37]
  wire  csignals_0 = _T_35 | _T_326; // @[Lookup.scala 33:37]
  wire [2:0] _T_327 = _T_229 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_328 = _T_227 ? 3'h5 : _T_327; // @[Lookup.scala 33:37]
  wire [2:0] _T_329 = _T_225 ? 3'h5 : _T_328; // @[Lookup.scala 33:37]
  wire [2:0] _T_330 = _T_223 ? 3'h5 : _T_329; // @[Lookup.scala 33:37]
  wire [2:0] _T_331 = _T_221 ? 3'h5 : _T_330; // @[Lookup.scala 33:37]
  wire [2:0] _T_332 = _T_219 ? 3'h5 : _T_331; // @[Lookup.scala 33:37]
  wire [2:0] _T_333 = _T_217 ? 3'h5 : _T_332; // @[Lookup.scala 33:37]
  wire [2:0] _T_334 = _T_215 ? 3'h5 : _T_333; // @[Lookup.scala 33:37]
  wire [2:0] _T_335 = _T_213 ? 3'h5 : _T_334; // @[Lookup.scala 33:37]
  wire [2:0] _T_336 = _T_211 ? 3'h5 : _T_335; // @[Lookup.scala 33:37]
  wire [2:0] _T_337 = _T_209 ? 3'h5 : _T_336; // @[Lookup.scala 33:37]
  wire [2:0] _T_338 = _T_207 ? 3'h5 : _T_337; // @[Lookup.scala 33:37]
  wire [2:0] _T_339 = _T_205 ? 3'h5 : _T_338; // @[Lookup.scala 33:37]
  wire [2:0] _T_340 = _T_203 ? 3'h5 : _T_339; // @[Lookup.scala 33:37]
  wire [2:0] _T_341 = _T_201 ? 3'h5 : _T_340; // @[Lookup.scala 33:37]
  wire [2:0] _T_342 = _T_199 ? 3'h5 : _T_341; // @[Lookup.scala 33:37]
  wire [2:0] _T_343 = _T_197 ? 3'h5 : _T_342; // @[Lookup.scala 33:37]
  wire [2:0] _T_344 = _T_195 ? 3'h5 : _T_343; // @[Lookup.scala 33:37]
  wire [2:0] _T_345 = _T_193 ? 3'h5 : _T_344; // @[Lookup.scala 33:37]
  wire [2:0] _T_346 = _T_191 ? 3'h5 : _T_345; // @[Lookup.scala 33:37]
  wire [2:0] _T_347 = _T_189 ? 3'h5 : _T_346; // @[Lookup.scala 33:37]
  wire [2:0] _T_348 = _T_187 ? 3'h5 : _T_347; // @[Lookup.scala 33:37]
  wire [2:0] _T_349 = _T_185 ? 3'h5 : _T_348; // @[Lookup.scala 33:37]
  wire [2:0] _T_350 = _T_183 ? 3'h5 : _T_349; // @[Lookup.scala 33:37]
  wire [2:0] _T_351 = _T_181 ? 3'h3 : _T_350; // @[Lookup.scala 33:37]
  wire [2:0] _T_352 = _T_179 ? 3'h3 : _T_351; // @[Lookup.scala 33:37]
  wire [2:0] _T_353 = _T_177 ? 3'h3 : _T_352; // @[Lookup.scala 33:37]
  wire [2:0] _T_354 = _T_175 ? 3'h3 : _T_353; // @[Lookup.scala 33:37]
  wire [2:0] _T_355 = _T_173 ? 3'h3 : _T_354; // @[Lookup.scala 33:37]
  wire [2:0] _T_356 = _T_171 ? 3'h3 : _T_355; // @[Lookup.scala 33:37]
  wire [2:0] _T_357 = _T_169 ? 3'h3 : _T_356; // @[Lookup.scala 33:37]
  wire [2:0] _T_358 = _T_167 ? 3'h3 : _T_357; // @[Lookup.scala 33:37]
  wire [2:0] _T_359 = _T_165 ? 3'h3 : _T_358; // @[Lookup.scala 33:37]
  wire [2:0] _T_360 = _T_163 ? 3'h3 : _T_359; // @[Lookup.scala 33:37]
  wire [2:0] _T_361 = _T_161 ? 3'h3 : _T_360; // @[Lookup.scala 33:37]
  wire [2:0] _T_362 = _T_159 ? 3'h3 : _T_361; // @[Lookup.scala 33:37]
  wire [2:0] _T_363 = _T_157 ? 3'h3 : _T_362; // @[Lookup.scala 33:37]
  wire [2:0] _T_364 = _T_155 ? 3'h3 : _T_363; // @[Lookup.scala 33:37]
  wire [2:0] _T_365 = _T_153 ? 3'h4 : _T_364; // @[Lookup.scala 33:37]
  wire [2:0] _T_366 = _T_151 ? 3'h4 : _T_365; // @[Lookup.scala 33:37]
  wire [2:0] _T_367 = _T_149 ? 3'h4 : _T_366; // @[Lookup.scala 33:37]
  wire [2:0] _T_368 = _T_147 ? 3'h4 : _T_367; // @[Lookup.scala 33:37]
  wire [2:0] _T_369 = _T_145 ? 3'h4 : _T_368; // @[Lookup.scala 33:37]
  wire [2:0] _T_370 = _T_143 ? 3'h4 : _T_369; // @[Lookup.scala 33:37]
  wire [2:0] _T_371 = _T_141 ? 3'h4 : _T_370; // @[Lookup.scala 33:37]
  wire [2:0] _T_372 = _T_139 ? 3'h4 : _T_371; // @[Lookup.scala 33:37]
  wire [2:0] _T_373 = _T_137 ? 3'h4 : _T_372; // @[Lookup.scala 33:37]
  wire [2:0] _T_374 = _T_135 ? 3'h4 : _T_373; // @[Lookup.scala 33:37]
  wire [2:0] _T_375 = _T_133 ? 3'h4 : _T_374; // @[Lookup.scala 33:37]
  wire [2:0] _T_376 = _T_131 ? 3'h4 : _T_375; // @[Lookup.scala 33:37]
  wire [2:0] _T_377 = _T_129 ? 3'h4 : _T_376; // @[Lookup.scala 33:37]
  wire [2:0] _T_378 = _T_127 ? 3'h2 : _T_377; // @[Lookup.scala 33:37]
  wire [2:0] _T_379 = _T_125 ? 3'h2 : _T_378; // @[Lookup.scala 33:37]
  wire [2:0] _T_380 = _T_123 ? 3'h2 : _T_379; // @[Lookup.scala 33:37]
  wire [2:0] _T_381 = _T_121 ? 3'h2 : _T_380; // @[Lookup.scala 33:37]
  wire [2:0] _T_382 = _T_119 ? 3'h2 : _T_381; // @[Lookup.scala 33:37]
  wire [2:0] _T_383 = _T_117 ? 3'h2 : _T_382; // @[Lookup.scala 33:37]
  wire [2:0] _T_384 = _T_115 ? 3'h2 : _T_383; // @[Lookup.scala 33:37]
  wire [2:0] _T_385 = _T_113 ? 3'h2 : _T_384; // @[Lookup.scala 33:37]
  wire [2:0] _T_386 = _T_111 ? 3'h2 : _T_385; // @[Lookup.scala 33:37]
  wire [2:0] _T_387 = _T_109 ? 3'h2 : _T_386; // @[Lookup.scala 33:37]
  wire [2:0] _T_388 = _T_107 ? 3'h2 : _T_387; // @[Lookup.scala 33:37]
  wire [2:0] _T_389 = _T_105 ? 3'h2 : _T_388; // @[Lookup.scala 33:37]
  wire [2:0] _T_390 = _T_103 ? 3'h1 : _T_389; // @[Lookup.scala 33:37]
  wire [2:0] _T_391 = _T_101 ? 3'h1 : _T_390; // @[Lookup.scala 33:37]
  wire [2:0] _T_392 = _T_99 ? 3'h1 : _T_391; // @[Lookup.scala 33:37]
  wire [2:0] _T_393 = _T_97 ? 3'h1 : _T_392; // @[Lookup.scala 33:37]
  wire [2:0] _T_394 = _T_95 ? 3'h1 : _T_393; // @[Lookup.scala 33:37]
  wire [2:0] _T_395 = _T_93 ? 3'h1 : _T_394; // @[Lookup.scala 33:37]
  wire [2:0] _T_396 = _T_91 ? 3'h1 : _T_395; // @[Lookup.scala 33:37]
  wire [2:0] _T_397 = _T_89 ? 3'h1 : _T_396; // @[Lookup.scala 33:37]
  wire [2:0] _T_398 = _T_87 ? 3'h1 : _T_397; // @[Lookup.scala 33:37]
  wire [2:0] _T_399 = _T_85 ? 3'h1 : _T_398; // @[Lookup.scala 33:37]
  wire [2:0] _T_400 = _T_83 ? 3'h1 : _T_399; // @[Lookup.scala 33:37]
  wire [2:0] _T_401 = _T_81 ? 3'h1 : _T_400; // @[Lookup.scala 33:37]
  wire [2:0] _T_402 = _T_79 ? 3'h1 : _T_401; // @[Lookup.scala 33:37]
  wire [2:0] _T_403 = _T_77 ? 3'h1 : _T_402; // @[Lookup.scala 33:37]
  wire [2:0] _T_404 = _T_75 ? 3'h1 : _T_403; // @[Lookup.scala 33:37]
  wire [2:0] _T_405 = _T_73 ? 3'h1 : _T_404; // @[Lookup.scala 33:37]
  wire [2:0] _T_406 = _T_71 ? 3'h1 : _T_405; // @[Lookup.scala 33:37]
  wire [2:0] _T_407 = _T_69 ? 3'h1 : _T_406; // @[Lookup.scala 33:37]
  wire [2:0] _T_408 = _T_67 ? 3'h1 : _T_407; // @[Lookup.scala 33:37]
  wire [2:0] _T_409 = _T_65 ? 3'h1 : _T_408; // @[Lookup.scala 33:37]
  wire [2:0] _T_410 = _T_63 ? 3'h1 : _T_409; // @[Lookup.scala 33:37]
  wire [2:0] _T_411 = _T_61 ? 3'h1 : _T_410; // @[Lookup.scala 33:37]
  wire [2:0] _T_412 = _T_59 ? 3'h1 : _T_411; // @[Lookup.scala 33:37]
  wire [2:0] _T_413 = _T_57 ? 3'h1 : _T_412; // @[Lookup.scala 33:37]
  wire [2:0] _T_414 = _T_55 ? 3'h1 : _T_413; // @[Lookup.scala 33:37]
  wire [2:0] _T_415 = _T_53 ? 3'h1 : _T_414; // @[Lookup.scala 33:37]
  wire [2:0] _T_416 = _T_51 ? 3'h1 : _T_415; // @[Lookup.scala 33:37]
  wire [2:0] _T_417 = _T_49 ? 3'h1 : _T_416; // @[Lookup.scala 33:37]
  wire [2:0] _T_418 = _T_47 ? 3'h1 : _T_417; // @[Lookup.scala 33:37]
  wire [2:0] _T_419 = _T_45 ? 3'h1 : _T_418; // @[Lookup.scala 33:37]
  wire [2:0] _T_420 = _T_43 ? 3'h1 : _T_419; // @[Lookup.scala 33:37]
  wire [2:0] _T_421 = _T_41 ? 3'h1 : _T_420; // @[Lookup.scala 33:37]
  wire [2:0] _T_422 = _T_39 ? 3'h1 : _T_421; // @[Lookup.scala 33:37]
  wire [2:0] _T_423 = _T_37 ? 3'h1 : _T_422; // @[Lookup.scala 33:37]
  wire [2:0] csignals_1 = _T_35 ? 3'h1 : _T_423; // @[Lookup.scala 33:37]
  wire [4:0] _T_424 = _T_229 ? 5'h18 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_425 = _T_227 ? 5'h17 : _T_424; // @[Lookup.scala 33:37]
  wire [4:0] _T_426 = _T_225 ? 5'h16 : _T_425; // @[Lookup.scala 33:37]
  wire [4:0] _T_427 = _T_223 ? 5'h15 : _T_426; // @[Lookup.scala 33:37]
  wire [4:0] _T_428 = _T_221 ? 5'h14 : _T_427; // @[Lookup.scala 33:37]
  wire [4:0] _T_429 = _T_219 ? 5'h13 : _T_428; // @[Lookup.scala 33:37]
  wire [4:0] _T_430 = _T_217 ? 5'h12 : _T_429; // @[Lookup.scala 33:37]
  wire [4:0] _T_431 = _T_215 ? 5'h11 : _T_430; // @[Lookup.scala 33:37]
  wire [4:0] _T_432 = _T_213 ? 5'h10 : _T_431; // @[Lookup.scala 33:37]
  wire [4:0] _T_433 = _T_211 ? 5'hf : _T_432; // @[Lookup.scala 33:37]
  wire [4:0] _T_434 = _T_209 ? 5'he : _T_433; // @[Lookup.scala 33:37]
  wire [4:0] _T_435 = _T_207 ? 5'hd : _T_434; // @[Lookup.scala 33:37]
  wire [4:0] _T_436 = _T_205 ? 5'h7 : _T_435; // @[Lookup.scala 33:37]
  wire [4:0] _T_437 = _T_203 ? 5'h6 : _T_436; // @[Lookup.scala 33:37]
  wire [4:0] _T_438 = _T_201 ? 5'h5 : _T_437; // @[Lookup.scala 33:37]
  wire [4:0] _T_439 = _T_199 ? 5'h8 : _T_438; // @[Lookup.scala 33:37]
  wire [4:0] _T_440 = _T_197 ? 5'hb : _T_439; // @[Lookup.scala 33:37]
  wire [4:0] _T_441 = _T_195 ? 5'hc : _T_440; // @[Lookup.scala 33:37]
  wire [4:0] _T_442 = _T_193 ? 5'ha : _T_441; // @[Lookup.scala 33:37]
  wire [4:0] _T_443 = _T_191 ? 5'h4 : _T_442; // @[Lookup.scala 33:37]
  wire [4:0] _T_444 = _T_189 ? 5'h3 : _T_443; // @[Lookup.scala 33:37]
  wire [4:0] _T_445 = _T_187 ? 5'h2 : _T_444; // @[Lookup.scala 33:37]
  wire [4:0] _T_446 = _T_185 ? 5'h9 : _T_445; // @[Lookup.scala 33:37]
  wire [4:0] _T_447 = _T_183 ? 5'h1 : _T_446; // @[Lookup.scala 33:37]
  wire [4:0] _T_448 = _T_181 ? 5'h1f : _T_447; // @[Lookup.scala 33:37]
  wire [4:0] _T_449 = _T_179 ? 5'h17 : _T_448; // @[Lookup.scala 33:37]
  wire [4:0] _T_450 = _T_177 ? 5'hf : _T_449; // @[Lookup.scala 33:37]
  wire [4:0] _T_451 = _T_175 ? 5'he : _T_450; // @[Lookup.scala 33:37]
  wire [4:0] _T_452 = _T_173 ? 5'h18 : _T_451; // @[Lookup.scala 33:37]
  wire [4:0] _T_453 = _T_171 ? 5'h1a : _T_452; // @[Lookup.scala 33:37]
  wire [4:0] _T_454 = _T_169 ? 5'h1e : _T_453; // @[Lookup.scala 33:37]
  wire [4:0] _T_455 = _T_167 ? 5'h7 : _T_454; // @[Lookup.scala 33:37]
  wire [4:0] _T_456 = _T_165 ? 5'h6 : _T_455; // @[Lookup.scala 33:37]
  wire [4:0] _T_457 = _T_163 ? 5'h11 : _T_456; // @[Lookup.scala 33:37]
  wire [4:0] _T_458 = _T_161 ? 5'h10 : _T_457; // @[Lookup.scala 33:37]
  wire [4:0] _T_459 = _T_159 ? 5'h13 : _T_458; // @[Lookup.scala 33:37]
  wire [4:0] _T_460 = _T_157 ? 5'h12 : _T_459; // @[Lookup.scala 33:37]
  wire [4:0] _T_461 = _T_155 ? 5'h16 : _T_460; // @[Lookup.scala 33:37]
  wire [4:0] _T_462 = _T_153 ? 5'h19 : _T_461; // @[Lookup.scala 33:37]
  wire [4:0] _T_463 = _T_151 ? 5'h17 : _T_462; // @[Lookup.scala 33:37]
  wire [4:0] _T_464 = _T_149 ? 5'h15 : _T_463; // @[Lookup.scala 33:37]
  wire [4:0] _T_465 = _T_147 ? 5'h13 : _T_464; // @[Lookup.scala 33:37]
  wire [4:0] _T_466 = _T_145 ? 5'h11 : _T_465; // @[Lookup.scala 33:37]
  wire [4:0] _T_467 = _T_143 ? 5'hf : _T_466; // @[Lookup.scala 33:37]
  wire [4:0] _T_468 = _T_141 ? 5'hd : _T_467; // @[Lookup.scala 33:37]
  wire [4:0] _T_469 = _T_139 ? 5'hb : _T_468; // @[Lookup.scala 33:37]
  wire [4:0] _T_470 = _T_137 ? 5'h8 : _T_469; // @[Lookup.scala 33:37]
  wire [4:0] _T_471 = _T_135 ? 5'h7 : _T_470; // @[Lookup.scala 33:37]
  wire [4:0] _T_472 = _T_133 ? 5'h5 : _T_471; // @[Lookup.scala 33:37]
  wire [4:0] _T_473 = _T_131 ? 5'h2 : _T_472; // @[Lookup.scala 33:37]
  wire [4:0] _T_474 = _T_129 ? 5'h0 : _T_473; // @[Lookup.scala 33:37]
  wire [4:0] _T_475 = _T_127 ? 5'hb : _T_474; // @[Lookup.scala 33:37]
  wire [4:0] _T_476 = _T_125 ? 5'ha : _T_475; // @[Lookup.scala 33:37]
  wire [4:0] _T_477 = _T_123 ? 5'h9 : _T_476; // @[Lookup.scala 33:37]
  wire [4:0] _T_478 = _T_121 ? 5'h8 : _T_477; // @[Lookup.scala 33:37]
  wire [4:0] _T_479 = _T_119 ? 5'h7 : _T_478; // @[Lookup.scala 33:37]
  wire [4:0] _T_480 = _T_117 ? 5'h6 : _T_479; // @[Lookup.scala 33:37]
  wire [4:0] _T_481 = _T_115 ? 5'h5 : _T_480; // @[Lookup.scala 33:37]
  wire [4:0] _T_482 = _T_113 ? 5'h4 : _T_481; // @[Lookup.scala 33:37]
  wire [4:0] _T_483 = _T_111 ? 5'h3 : _T_482; // @[Lookup.scala 33:37]
  wire [4:0] _T_484 = _T_109 ? 5'h2 : _T_483; // @[Lookup.scala 33:37]
  wire [4:0] _T_485 = _T_107 ? 5'h1 : _T_484; // @[Lookup.scala 33:37]
  wire [4:0] _T_486 = _T_105 ? 5'h0 : _T_485; // @[Lookup.scala 33:37]
  wire [4:0] _T_487 = _T_103 ? 5'h17 : _T_486; // @[Lookup.scala 33:37]
  wire [4:0] _T_488 = _T_101 ? 5'h17 : _T_487; // @[Lookup.scala 33:37]
  wire [4:0] _T_489 = _T_99 ? 5'h16 : _T_488; // @[Lookup.scala 33:37]
  wire [4:0] _T_490 = _T_97 ? 5'h15 : _T_489; // @[Lookup.scala 33:37]
  wire [4:0] _T_491 = _T_95 ? 5'h14 : _T_490; // @[Lookup.scala 33:37]
  wire [4:0] _T_492 = _T_93 ? 5'h13 : _T_491; // @[Lookup.scala 33:37]
  wire [4:0] _T_493 = _T_91 ? 5'h12 : _T_492; // @[Lookup.scala 33:37]
  wire [4:0] _T_494 = _T_89 ? 5'h11 : _T_493; // @[Lookup.scala 33:37]
  wire [4:0] _T_495 = _T_87 ? 5'h10 : _T_494; // @[Lookup.scala 33:37]
  wire [4:0] _T_496 = _T_85 ? 5'hd : _T_495; // @[Lookup.scala 33:37]
  wire [4:0] _T_497 = _T_83 ? 5'hc : _T_496; // @[Lookup.scala 33:37]
  wire [4:0] _T_498 = _T_81 ? 5'h7 : _T_497; // @[Lookup.scala 33:37]
  wire [4:0] _T_499 = _T_79 ? 5'h6 : _T_498; // @[Lookup.scala 33:37]
  wire [4:0] _T_500 = _T_77 ? 5'h5 : _T_499; // @[Lookup.scala 33:37]
  wire [4:0] _T_501 = _T_75 ? 5'h0 : _T_500; // @[Lookup.scala 33:37]
  wire [4:0] _T_502 = _T_73 ? 5'he : _T_501; // @[Lookup.scala 33:37]
  wire [4:0] _T_503 = _T_71 ? 5'h2 : _T_502; // @[Lookup.scala 33:37]
  wire [4:0] _T_504 = _T_69 ? 5'h3 : _T_503; // @[Lookup.scala 33:37]
  wire [4:0] _T_505 = _T_67 ? 5'h4 : _T_504; // @[Lookup.scala 33:37]
  wire [4:0] _T_506 = _T_65 ? 5'h3 : _T_505; // @[Lookup.scala 33:37]
  wire [4:0] _T_507 = _T_63 ? 5'h4 : _T_506; // @[Lookup.scala 33:37]
  wire [4:0] _T_508 = _T_61 ? 5'h2 : _T_507; // @[Lookup.scala 33:37]
  wire [4:0] _T_509 = _T_59 ? 5'ha : _T_508; // @[Lookup.scala 33:37]
  wire [4:0] _T_510 = _T_57 ? 5'h9 : _T_509; // @[Lookup.scala 33:37]
  wire [4:0] _T_511 = _T_55 ? 5'h8 : _T_510; // @[Lookup.scala 33:37]
  wire [4:0] _T_512 = _T_53 ? 5'h7 : _T_511; // @[Lookup.scala 33:37]
  wire [4:0] _T_513 = _T_51 ? 5'h6 : _T_512; // @[Lookup.scala 33:37]
  wire [4:0] _T_514 = _T_49 ? 5'h5 : _T_513; // @[Lookup.scala 33:37]
  wire [4:0] _T_515 = _T_47 ? 5'ha : _T_514; // @[Lookup.scala 33:37]
  wire [4:0] _T_516 = _T_45 ? 5'h9 : _T_515; // @[Lookup.scala 33:37]
  wire [4:0] _T_517 = _T_43 ? 5'h1 : _T_516; // @[Lookup.scala 33:37]
  wire [4:0] _T_518 = _T_41 ? 5'hf : _T_517; // @[Lookup.scala 33:37]
  wire [4:0] _T_519 = _T_39 ? 5'h0 : _T_518; // @[Lookup.scala 33:37]
  wire [4:0] _T_520 = _T_37 ? 5'he : _T_519; // @[Lookup.scala 33:37]
  wire [4:0] csignals_2 = _T_35 ? 5'hb : _T_520; // @[Lookup.scala 33:37]
  wire [1:0] _T_521 = _T_229 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_522 = _T_227 ? 2'h1 : _T_521; // @[Lookup.scala 33:37]
  wire [1:0] _T_523 = _T_225 ? 2'h1 : _T_522; // @[Lookup.scala 33:37]
  wire [1:0] _T_524 = _T_223 ? 2'h1 : _T_523; // @[Lookup.scala 33:37]
  wire [1:0] _T_525 = _T_221 ? 2'h1 : _T_524; // @[Lookup.scala 33:37]
  wire [1:0] _T_526 = _T_219 ? 2'h1 : _T_525; // @[Lookup.scala 33:37]
  wire [1:0] _T_527 = _T_217 ? 2'h1 : _T_526; // @[Lookup.scala 33:37]
  wire [1:0] _T_528 = _T_215 ? 2'h1 : _T_527; // @[Lookup.scala 33:37]
  wire [1:0] _T_529 = _T_213 ? 2'h1 : _T_528; // @[Lookup.scala 33:37]
  wire [1:0] _T_530 = _T_211 ? 2'h1 : _T_529; // @[Lookup.scala 33:37]
  wire [1:0] _T_531 = _T_209 ? 2'h1 : _T_530; // @[Lookup.scala 33:37]
  wire [1:0] _T_532 = _T_207 ? 2'h1 : _T_531; // @[Lookup.scala 33:37]
  wire [1:0] _T_533 = _T_205 ? 2'h0 : _T_532; // @[Lookup.scala 33:37]
  wire [1:0] _T_534 = _T_203 ? 2'h0 : _T_533; // @[Lookup.scala 33:37]
  wire [1:0] _T_535 = _T_201 ? 2'h0 : _T_534; // @[Lookup.scala 33:37]
  wire [1:0] _T_536 = _T_199 ? 2'h0 : _T_535; // @[Lookup.scala 33:37]
  wire [1:0] _T_537 = _T_197 ? 2'h0 : _T_536; // @[Lookup.scala 33:37]
  wire [1:0] _T_538 = _T_195 ? 2'h0 : _T_537; // @[Lookup.scala 33:37]
  wire [1:0] _T_539 = _T_193 ? 2'h3 : _T_538; // @[Lookup.scala 33:37]
  wire [1:0] _T_540 = _T_191 ? 2'h2 : _T_539; // @[Lookup.scala 33:37]
  wire [1:0] _T_541 = _T_189 ? 2'h0 : _T_540; // @[Lookup.scala 33:37]
  wire [1:0] _T_542 = _T_187 ? 2'h0 : _T_541; // @[Lookup.scala 33:37]
  wire [1:0] _T_543 = _T_185 ? 2'h0 : _T_542; // @[Lookup.scala 33:37]
  wire [1:0] _T_544 = _T_183 ? 2'h0 : _T_543; // @[Lookup.scala 33:37]
  wire [1:0] _T_545 = _T_181 ? 2'h3 : _T_544; // @[Lookup.scala 33:37]
  wire [1:0] _T_546 = _T_179 ? 2'h3 : _T_545; // @[Lookup.scala 33:37]
  wire [1:0] _T_547 = _T_177 ? 2'h3 : _T_546; // @[Lookup.scala 33:37]
  wire [1:0] _T_548 = _T_175 ? 2'h3 : _T_547; // @[Lookup.scala 33:37]
  wire [1:0] _T_549 = _T_173 ? 2'h3 : _T_548; // @[Lookup.scala 33:37]
  wire [1:0] _T_550 = _T_171 ? 2'h3 : _T_549; // @[Lookup.scala 33:37]
  wire [1:0] _T_551 = _T_169 ? 2'h3 : _T_550; // @[Lookup.scala 33:37]
  wire [1:0] _T_552 = _T_167 ? 2'h3 : _T_551; // @[Lookup.scala 33:37]
  wire [1:0] _T_553 = _T_165 ? 2'h3 : _T_552; // @[Lookup.scala 33:37]
  wire [1:0] _T_554 = _T_163 ? 2'h3 : _T_553; // @[Lookup.scala 33:37]
  wire [1:0] _T_555 = _T_161 ? 2'h3 : _T_554; // @[Lookup.scala 33:37]
  wire [1:0] _T_556 = _T_159 ? 2'h3 : _T_555; // @[Lookup.scala 33:37]
  wire [1:0] _T_557 = _T_157 ? 2'h3 : _T_556; // @[Lookup.scala 33:37]
  wire [1:0] _T_558 = _T_155 ? 2'h3 : _T_557; // @[Lookup.scala 33:37]
  wire [1:0] _T_559 = _T_153 ? 2'h1 : _T_558; // @[Lookup.scala 33:37]
  wire [1:0] _T_560 = _T_151 ? 2'h1 : _T_559; // @[Lookup.scala 33:37]
  wire [1:0] _T_561 = _T_149 ? 2'h1 : _T_560; // @[Lookup.scala 33:37]
  wire [1:0] _T_562 = _T_147 ? 2'h1 : _T_561; // @[Lookup.scala 33:37]
  wire [1:0] _T_563 = _T_145 ? 2'h1 : _T_562; // @[Lookup.scala 33:37]
  wire [1:0] _T_564 = _T_143 ? 2'h1 : _T_563; // @[Lookup.scala 33:37]
  wire [1:0] _T_565 = _T_141 ? 2'h1 : _T_564; // @[Lookup.scala 33:37]
  wire [1:0] _T_566 = _T_139 ? 2'h1 : _T_565; // @[Lookup.scala 33:37]
  wire [1:0] _T_567 = _T_137 ? 2'h1 : _T_566; // @[Lookup.scala 33:37]
  wire [1:0] _T_568 = _T_135 ? 2'h1 : _T_567; // @[Lookup.scala 33:37]
  wire [1:0] _T_569 = _T_133 ? 2'h1 : _T_568; // @[Lookup.scala 33:37]
  wire [1:0] _T_570 = _T_131 ? 2'h0 : _T_569; // @[Lookup.scala 33:37]
  wire [1:0] _T_571 = _T_129 ? 2'h0 : _T_570; // @[Lookup.scala 33:37]
  wire [1:0] _T_572 = _T_127 ? 2'h1 : _T_571; // @[Lookup.scala 33:37]
  wire [1:0] _T_573 = _T_125 ? 2'h1 : _T_572; // @[Lookup.scala 33:37]
  wire [1:0] _T_574 = _T_123 ? 2'h1 : _T_573; // @[Lookup.scala 33:37]
  wire [1:0] _T_575 = _T_121 ? 2'h1 : _T_574; // @[Lookup.scala 33:37]
  wire [1:0] _T_576 = _T_119 ? 2'h1 : _T_575; // @[Lookup.scala 33:37]
  wire [1:0] _T_577 = _T_117 ? 2'h1 : _T_576; // @[Lookup.scala 33:37]
  wire [1:0] _T_578 = _T_115 ? 2'h1 : _T_577; // @[Lookup.scala 33:37]
  wire [1:0] _T_579 = _T_113 ? 2'h1 : _T_578; // @[Lookup.scala 33:37]
  wire [1:0] _T_580 = _T_111 ? 2'h1 : _T_579; // @[Lookup.scala 33:37]
  wire [1:0] _T_581 = _T_109 ? 2'h1 : _T_580; // @[Lookup.scala 33:37]
  wire [1:0] _T_582 = _T_107 ? 2'h1 : _T_581; // @[Lookup.scala 33:37]
  wire [1:0] _T_583 = _T_105 ? 2'h1 : _T_582; // @[Lookup.scala 33:37]
  wire [1:0] _T_584 = _T_103 ? 2'h2 : _T_583; // @[Lookup.scala 33:37]
  wire [1:0] _T_585 = _T_101 ? 2'h2 : _T_584; // @[Lookup.scala 33:37]
  wire [1:0] _T_586 = _T_99 ? 2'h1 : _T_585; // @[Lookup.scala 33:37]
  wire [1:0] _T_587 = _T_97 ? 2'h1 : _T_586; // @[Lookup.scala 33:37]
  wire [1:0] _T_588 = _T_95 ? 2'h2 : _T_587; // @[Lookup.scala 33:37]
  wire [1:0] _T_589 = _T_93 ? 2'h2 : _T_588; // @[Lookup.scala 33:37]
  wire [1:0] _T_590 = _T_91 ? 2'h2 : _T_589; // @[Lookup.scala 33:37]
  wire [1:0] _T_591 = _T_89 ? 2'h1 : _T_590; // @[Lookup.scala 33:37]
  wire [1:0] _T_592 = _T_87 ? 2'h1 : _T_591; // @[Lookup.scala 33:37]
  wire [1:0] _T_593 = _T_85 ? 2'h1 : _T_592; // @[Lookup.scala 33:37]
  wire [1:0] _T_594 = _T_83 ? 2'h1 : _T_593; // @[Lookup.scala 33:37]
  wire [1:0] _T_595 = _T_81 ? 2'h1 : _T_594; // @[Lookup.scala 33:37]
  wire [1:0] _T_596 = _T_79 ? 2'h1 : _T_595; // @[Lookup.scala 33:37]
  wire [1:0] _T_597 = _T_77 ? 2'h1 : _T_596; // @[Lookup.scala 33:37]
  wire [1:0] _T_598 = _T_75 ? 2'h1 : _T_597; // @[Lookup.scala 33:37]
  wire [1:0] _T_599 = _T_73 ? 2'h1 : _T_598; // @[Lookup.scala 33:37]
  wire [1:0] _T_600 = _T_71 ? 2'h2 : _T_599; // @[Lookup.scala 33:37]
  wire [1:0] _T_601 = _T_69 ? 2'h2 : _T_600; // @[Lookup.scala 33:37]
  wire [1:0] _T_602 = _T_67 ? 2'h2 : _T_601; // @[Lookup.scala 33:37]
  wire [1:0] _T_603 = _T_65 ? 2'h2 : _T_602; // @[Lookup.scala 33:37]
  wire [1:0] _T_604 = _T_63 ? 2'h2 : _T_603; // @[Lookup.scala 33:37]
  wire [1:0] _T_605 = _T_61 ? 2'h2 : _T_604; // @[Lookup.scala 33:37]
  wire [1:0] _T_606 = _T_59 ? 2'h1 : _T_605; // @[Lookup.scala 33:37]
  wire [1:0] _T_607 = _T_57 ? 2'h1 : _T_606; // @[Lookup.scala 33:37]
  wire [1:0] _T_608 = _T_55 ? 2'h1 : _T_607; // @[Lookup.scala 33:37]
  wire [1:0] _T_609 = _T_53 ? 2'h1 : _T_608; // @[Lookup.scala 33:37]
  wire [1:0] _T_610 = _T_51 ? 2'h1 : _T_609; // @[Lookup.scala 33:37]
  wire [1:0] _T_611 = _T_49 ? 2'h1 : _T_610; // @[Lookup.scala 33:37]
  wire [1:0] _T_612 = _T_47 ? 2'h1 : _T_611; // @[Lookup.scala 33:37]
  wire [1:0] _T_613 = _T_45 ? 2'h1 : _T_612; // @[Lookup.scala 33:37]
  wire [1:0] _T_614 = _T_43 ? 2'h1 : _T_613; // @[Lookup.scala 33:37]
  wire [1:0] _T_615 = _T_41 ? 2'h1 : _T_614; // @[Lookup.scala 33:37]
  wire [1:0] _T_616 = _T_39 ? 2'h1 : _T_615; // @[Lookup.scala 33:37]
  wire [1:0] _T_617 = _T_37 ? 2'h1 : _T_616; // @[Lookup.scala 33:37]
  wire [1:0] csignals_3 = _T_35 ? 2'h0 : _T_617; // @[Lookup.scala 33:37]
  wire [2:0] _T_618 = _T_229 ? 3'h3 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_619 = _T_227 ? 3'h3 : _T_618; // @[Lookup.scala 33:37]
  wire [2:0] _T_620 = _T_225 ? 3'h3 : _T_619; // @[Lookup.scala 33:37]
  wire [2:0] _T_621 = _T_223 ? 3'h3 : _T_620; // @[Lookup.scala 33:37]
  wire [2:0] _T_622 = _T_221 ? 3'h3 : _T_621; // @[Lookup.scala 33:37]
  wire [2:0] _T_623 = _T_219 ? 3'h3 : _T_622; // @[Lookup.scala 33:37]
  wire [2:0] _T_624 = _T_217 ? 3'h2 : _T_623; // @[Lookup.scala 33:37]
  wire [2:0] _T_625 = _T_215 ? 3'h2 : _T_624; // @[Lookup.scala 33:37]
  wire [2:0] _T_626 = _T_213 ? 3'h2 : _T_625; // @[Lookup.scala 33:37]
  wire [2:0] _T_627 = _T_211 ? 3'h2 : _T_626; // @[Lookup.scala 33:37]
  wire [2:0] _T_628 = _T_209 ? 3'h2 : _T_627; // @[Lookup.scala 33:37]
  wire [2:0] _T_629 = _T_207 ? 3'h2 : _T_628; // @[Lookup.scala 33:37]
  wire [2:0] _T_630 = _T_205 ? 3'h0 : _T_629; // @[Lookup.scala 33:37]
  wire [2:0] _T_631 = _T_203 ? 3'h0 : _T_630; // @[Lookup.scala 33:37]
  wire [2:0] _T_632 = _T_201 ? 3'h0 : _T_631; // @[Lookup.scala 33:37]
  wire [2:0] _T_633 = _T_199 ? 3'h0 : _T_632; // @[Lookup.scala 33:37]
  wire [2:0] _T_634 = _T_197 ? 3'h0 : _T_633; // @[Lookup.scala 33:37]
  wire [2:0] _T_635 = _T_195 ? 3'h0 : _T_634; // @[Lookup.scala 33:37]
  wire [2:0] _T_636 = _T_193 ? 3'h7 : _T_635; // @[Lookup.scala 33:37]
  wire [2:0] _T_637 = _T_191 ? 3'h0 : _T_636; // @[Lookup.scala 33:37]
  wire [2:0] _T_638 = _T_189 ? 3'h0 : _T_637; // @[Lookup.scala 33:37]
  wire [2:0] _T_639 = _T_187 ? 3'h0 : _T_638; // @[Lookup.scala 33:37]
  wire [2:0] _T_640 = _T_185 ? 3'h0 : _T_639; // @[Lookup.scala 33:37]
  wire [2:0] _T_641 = _T_183 ? 3'h0 : _T_640; // @[Lookup.scala 33:37]
  wire [2:0] _T_642 = _T_181 ? 3'h2 : _T_641; // @[Lookup.scala 33:37]
  wire [2:0] _T_643 = _T_179 ? 3'h0 : _T_642; // @[Lookup.scala 33:37]
  wire [2:0] _T_644 = _T_177 ? 3'h2 : _T_643; // @[Lookup.scala 33:37]
  wire [2:0] _T_645 = _T_175 ? 3'h2 : _T_644; // @[Lookup.scala 33:37]
  wire [2:0] _T_646 = _T_173 ? 3'h2 : _T_645; // @[Lookup.scala 33:37]
  wire [2:0] _T_647 = _T_171 ? 3'h2 : _T_646; // @[Lookup.scala 33:37]
  wire [2:0] _T_648 = _T_169 ? 3'h2 : _T_647; // @[Lookup.scala 33:37]
  wire [2:0] _T_649 = _T_167 ? 3'h2 : _T_648; // @[Lookup.scala 33:37]
  wire [2:0] _T_650 = _T_165 ? 3'h2 : _T_649; // @[Lookup.scala 33:37]
  wire [2:0] _T_651 = _T_163 ? 3'h0 : _T_650; // @[Lookup.scala 33:37]
  wire [2:0] _T_652 = _T_161 ? 3'h0 : _T_651; // @[Lookup.scala 33:37]
  wire [2:0] _T_653 = _T_159 ? 3'h0 : _T_652; // @[Lookup.scala 33:37]
  wire [2:0] _T_654 = _T_157 ? 3'h0 : _T_653; // @[Lookup.scala 33:37]
  wire [2:0] _T_655 = _T_155 ? 3'h0 : _T_654; // @[Lookup.scala 33:37]
  wire [2:0] _T_656 = _T_153 ? 3'h2 : _T_655; // @[Lookup.scala 33:37]
  wire [2:0] _T_657 = _T_151 ? 3'h2 : _T_656; // @[Lookup.scala 33:37]
  wire [2:0] _T_658 = _T_149 ? 3'h2 : _T_657; // @[Lookup.scala 33:37]
  wire [2:0] _T_659 = _T_147 ? 3'h2 : _T_658; // @[Lookup.scala 33:37]
  wire [2:0] _T_660 = _T_145 ? 3'h2 : _T_659; // @[Lookup.scala 33:37]
  wire [2:0] _T_661 = _T_143 ? 3'h2 : _T_660; // @[Lookup.scala 33:37]
  wire [2:0] _T_662 = _T_141 ? 3'h2 : _T_661; // @[Lookup.scala 33:37]
  wire [2:0] _T_663 = _T_139 ? 3'h2 : _T_662; // @[Lookup.scala 33:37]
  wire [2:0] _T_664 = _T_137 ? 3'h2 : _T_663; // @[Lookup.scala 33:37]
  wire [2:0] _T_665 = _T_135 ? 3'h0 : _T_664; // @[Lookup.scala 33:37]
  wire [2:0] _T_666 = _T_133 ? 3'h0 : _T_665; // @[Lookup.scala 33:37]
  wire [2:0] _T_667 = _T_131 ? 3'h0 : _T_666; // @[Lookup.scala 33:37]
  wire [2:0] _T_668 = _T_129 ? 3'h0 : _T_667; // @[Lookup.scala 33:37]
  wire [2:0] _T_669 = _T_127 ? 3'h0 : _T_668; // @[Lookup.scala 33:37]
  wire [2:0] _T_670 = _T_125 ? 3'h0 : _T_669; // @[Lookup.scala 33:37]
  wire [2:0] _T_671 = _T_123 ? 3'h0 : _T_670; // @[Lookup.scala 33:37]
  wire [2:0] _T_672 = _T_121 ? 3'h0 : _T_671; // @[Lookup.scala 33:37]
  wire [2:0] _T_673 = _T_119 ? 3'h0 : _T_672; // @[Lookup.scala 33:37]
  wire [2:0] _T_674 = _T_117 ? 3'h0 : _T_673; // @[Lookup.scala 33:37]
  wire [2:0] _T_675 = _T_115 ? 3'h0 : _T_674; // @[Lookup.scala 33:37]
  wire [2:0] _T_676 = _T_113 ? 3'h0 : _T_675; // @[Lookup.scala 33:37]
  wire [2:0] _T_677 = _T_111 ? 3'h0 : _T_676; // @[Lookup.scala 33:37]
  wire [2:0] _T_678 = _T_109 ? 3'h0 : _T_677; // @[Lookup.scala 33:37]
  wire [2:0] _T_679 = _T_107 ? 3'h2 : _T_678; // @[Lookup.scala 33:37]
  wire [2:0] _T_680 = _T_105 ? 3'h2 : _T_679; // @[Lookup.scala 33:37]
  wire [2:0] _T_681 = _T_103 ? 3'h1 : _T_680; // @[Lookup.scala 33:37]
  wire [2:0] _T_682 = _T_101 ? 3'h6 : _T_681; // @[Lookup.scala 33:37]
  wire [2:0] _T_683 = _T_99 ? 3'h0 : _T_682; // @[Lookup.scala 33:37]
  wire [2:0] _T_684 = _T_97 ? 3'h2 : _T_683; // @[Lookup.scala 33:37]
  wire [2:0] _T_685 = _T_95 ? 3'h0 : _T_684; // @[Lookup.scala 33:37]
  wire [2:0] _T_686 = _T_93 ? 3'h0 : _T_685; // @[Lookup.scala 33:37]
  wire [2:0] _T_687 = _T_91 ? 3'h0 : _T_686; // @[Lookup.scala 33:37]
  wire [2:0] _T_688 = _T_89 ? 3'h0 : _T_687; // @[Lookup.scala 33:37]
  wire [2:0] _T_689 = _T_87 ? 3'h0 : _T_688; // @[Lookup.scala 33:37]
  wire [2:0] _T_690 = _T_85 ? 3'h2 : _T_689; // @[Lookup.scala 33:37]
  wire [2:0] _T_691 = _T_83 ? 3'h2 : _T_690; // @[Lookup.scala 33:37]
  wire [2:0] _T_692 = _T_81 ? 3'h5 : _T_691; // @[Lookup.scala 33:37]
  wire [2:0] _T_693 = _T_79 ? 3'h5 : _T_692; // @[Lookup.scala 33:37]
  wire [2:0] _T_694 = _T_77 ? 3'h5 : _T_693; // @[Lookup.scala 33:37]
  wire [2:0] _T_695 = _T_75 ? 3'h3 : _T_694; // @[Lookup.scala 33:37]
  wire [2:0] _T_696 = _T_73 ? 3'h3 : _T_695; // @[Lookup.scala 33:37]
  wire [2:0] _T_697 = _T_71 ? 3'h1 : _T_696; // @[Lookup.scala 33:37]
  wire [2:0] _T_698 = _T_69 ? 3'h1 : _T_697; // @[Lookup.scala 33:37]
  wire [2:0] _T_699 = _T_67 ? 3'h1 : _T_698; // @[Lookup.scala 33:37]
  wire [2:0] _T_700 = _T_65 ? 3'h6 : _T_699; // @[Lookup.scala 33:37]
  wire [2:0] _T_701 = _T_63 ? 3'h6 : _T_700; // @[Lookup.scala 33:37]
  wire [2:0] _T_702 = _T_61 ? 3'h6 : _T_701; // @[Lookup.scala 33:37]
  wire [2:0] _T_703 = _T_59 ? 3'h3 : _T_702; // @[Lookup.scala 33:37]
  wire [2:0] _T_704 = _T_57 ? 3'h3 : _T_703; // @[Lookup.scala 33:37]
  wire [2:0] _T_705 = _T_55 ? 3'h2 : _T_704; // @[Lookup.scala 33:37]
  wire [2:0] _T_706 = _T_53 ? 3'h2 : _T_705; // @[Lookup.scala 33:37]
  wire [2:0] _T_707 = _T_51 ? 3'h2 : _T_706; // @[Lookup.scala 33:37]
  wire [2:0] _T_708 = _T_49 ? 3'h2 : _T_707; // @[Lookup.scala 33:37]
  wire [2:0] _T_709 = _T_47 ? 3'h2 : _T_708; // @[Lookup.scala 33:37]
  wire [2:0] _T_710 = _T_45 ? 3'h2 : _T_709; // @[Lookup.scala 33:37]
  wire [2:0] _T_711 = _T_43 ? 3'h2 : _T_710; // @[Lookup.scala 33:37]
  wire [2:0] _T_712 = _T_41 ? 3'h2 : _T_711; // @[Lookup.scala 33:37]
  wire [2:0] _T_713 = _T_39 ? 3'h2 : _T_712; // @[Lookup.scala 33:37]
  wire [2:0] _T_714 = _T_37 ? 3'h2 : _T_713; // @[Lookup.scala 33:37]
  wire [2:0] csignals_4 = _T_35 ? 3'h4 : _T_714; // @[Lookup.scala 33:37]
  wire [1:0] _T_735 = _T_189 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_736 = _T_187 ? 2'h0 : _T_735; // @[Lookup.scala 33:37]
  wire [1:0] _T_737 = _T_185 ? 2'h0 : _T_736; // @[Lookup.scala 33:37]
  wire [1:0] _T_738 = _T_183 ? 2'h0 : _T_737; // @[Lookup.scala 33:37]
  wire [1:0] _T_739 = _T_181 ? 2'h2 : _T_738; // @[Lookup.scala 33:37]
  wire [1:0] _T_740 = _T_179 ? 2'h2 : _T_739; // @[Lookup.scala 33:37]
  wire [1:0] _T_741 = _T_177 ? 2'h0 : _T_740; // @[Lookup.scala 33:37]
  wire [1:0] _T_742 = _T_175 ? 2'h0 : _T_741; // @[Lookup.scala 33:37]
  wire [1:0] _T_743 = _T_173 ? 2'h0 : _T_742; // @[Lookup.scala 33:37]
  wire [1:0] _T_744 = _T_171 ? 2'h0 : _T_743; // @[Lookup.scala 33:37]
  wire [1:0] _T_745 = _T_169 ? 2'h0 : _T_744; // @[Lookup.scala 33:37]
  wire [1:0] _T_746 = _T_167 ? 2'h2 : _T_745; // @[Lookup.scala 33:37]
  wire [1:0] _T_747 = _T_165 ? 2'h2 : _T_746; // @[Lookup.scala 33:37]
  wire [1:0] _T_748 = _T_163 ? 2'h2 : _T_747; // @[Lookup.scala 33:37]
  wire [1:0] _T_749 = _T_161 ? 2'h2 : _T_748; // @[Lookup.scala 33:37]
  wire [1:0] _T_750 = _T_159 ? 2'h2 : _T_749; // @[Lookup.scala 33:37]
  wire [1:0] _T_751 = _T_157 ? 2'h2 : _T_750; // @[Lookup.scala 33:37]
  wire [1:0] _T_752 = _T_155 ? 2'h2 : _T_751; // @[Lookup.scala 33:37]
  wire [1:0] _T_753 = _T_153 ? 2'h0 : _T_752; // @[Lookup.scala 33:37]
  wire [1:0] _T_754 = _T_151 ? 2'h0 : _T_753; // @[Lookup.scala 33:37]
  wire [1:0] _T_755 = _T_149 ? 2'h0 : _T_754; // @[Lookup.scala 33:37]
  wire [1:0] _T_756 = _T_147 ? 2'h0 : _T_755; // @[Lookup.scala 33:37]
  wire [1:0] _T_757 = _T_145 ? 2'h0 : _T_756; // @[Lookup.scala 33:37]
  wire [1:0] _T_758 = _T_143 ? 2'h0 : _T_757; // @[Lookup.scala 33:37]
  wire [1:0] _T_759 = _T_141 ? 2'h0 : _T_758; // @[Lookup.scala 33:37]
  wire [1:0] _T_760 = _T_139 ? 2'h0 : _T_759; // @[Lookup.scala 33:37]
  wire [1:0] _T_761 = _T_137 ? 2'h1 : _T_760; // @[Lookup.scala 33:37]
  wire [1:0] _T_762 = _T_135 ? 2'h0 : _T_761; // @[Lookup.scala 33:37]
  wire [1:0] _T_763 = _T_133 ? 2'h0 : _T_762; // @[Lookup.scala 33:37]
  wire [1:0] _T_764 = _T_131 ? 2'h1 : _T_763; // @[Lookup.scala 33:37]
  wire [1:0] _T_765 = _T_129 ? 2'h1 : _T_764; // @[Lookup.scala 33:37]
  wire [1:0] _T_766 = _T_127 ? 2'h1 : _T_765; // @[Lookup.scala 33:37]
  wire [1:0] _T_767 = _T_125 ? 2'h0 : _T_766; // @[Lookup.scala 33:37]
  wire [1:0] _T_768 = _T_123 ? 2'h3 : _T_767; // @[Lookup.scala 33:37]
  wire [1:0] _T_769 = _T_121 ? 2'h0 : _T_768; // @[Lookup.scala 33:37]
  wire [1:0] _T_770 = _T_119 ? 2'h3 : _T_769; // @[Lookup.scala 33:37]
  wire [1:0] _T_771 = _T_117 ? 2'h3 : _T_770; // @[Lookup.scala 33:37]
  wire [1:0] _T_772 = _T_115 ? 2'h0 : _T_771; // @[Lookup.scala 33:37]
  wire [1:0] _T_773 = _T_113 ? 2'h0 : _T_772; // @[Lookup.scala 33:37]
  wire [1:0] _T_774 = _T_111 ? 2'h0 : _T_773; // @[Lookup.scala 33:37]
  wire [1:0] _T_775 = _T_109 ? 2'h0 : _T_774; // @[Lookup.scala 33:37]
  wire [1:0] _T_776 = _T_107 ? 2'h0 : _T_775; // @[Lookup.scala 33:37]
  wire [1:0] _T_777 = _T_105 ? 2'h0 : _T_776; // @[Lookup.scala 33:37]
  wire [1:0] _T_778 = _T_103 ? 2'h1 : _T_777; // @[Lookup.scala 33:37]
  wire [1:0] _T_779 = _T_101 ? 2'h1 : _T_778; // @[Lookup.scala 33:37]
  wire [1:0] _T_780 = _T_99 ? 2'h2 : _T_779; // @[Lookup.scala 33:37]
  wire [1:0] _T_781 = _T_97 ? 2'h2 : _T_780; // @[Lookup.scala 33:37]
  wire [1:0] _T_782 = _T_95 ? 2'h1 : _T_781; // @[Lookup.scala 33:37]
  wire [1:0] _T_783 = _T_93 ? 2'h1 : _T_782; // @[Lookup.scala 33:37]
  wire [1:0] _T_784 = _T_91 ? 2'h1 : _T_783; // @[Lookup.scala 33:37]
  wire [1:0] _T_785 = _T_89 ? 2'h1 : _T_784; // @[Lookup.scala 33:37]
  wire [1:0] _T_786 = _T_87 ? 2'h1 : _T_785; // @[Lookup.scala 33:37]
  wire [1:0] _T_787 = _T_85 ? 2'h1 : _T_786; // @[Lookup.scala 33:37]
  wire [1:0] _T_788 = _T_83 ? 2'h1 : _T_787; // @[Lookup.scala 33:37]
  wire [1:0] _T_789 = _T_81 ? 2'h2 : _T_788; // @[Lookup.scala 33:37]
  wire [1:0] _T_790 = _T_79 ? 2'h2 : _T_789; // @[Lookup.scala 33:37]
  wire [1:0] _T_791 = _T_77 ? 2'h2 : _T_790; // @[Lookup.scala 33:37]
  wire [1:0] _T_792 = _T_75 ? 2'h2 : _T_791; // @[Lookup.scala 33:37]
  wire [1:0] _T_793 = _T_73 ? 2'h2 : _T_792; // @[Lookup.scala 33:37]
  wire [1:0] _T_794 = _T_71 ? 2'h1 : _T_793; // @[Lookup.scala 33:37]
  wire [1:0] _T_795 = _T_69 ? 2'h1 : _T_794; // @[Lookup.scala 33:37]
  wire [1:0] _T_796 = _T_67 ? 2'h1 : _T_795; // @[Lookup.scala 33:37]
  wire [1:0] _T_797 = _T_65 ? 2'h1 : _T_796; // @[Lookup.scala 33:37]
  wire [1:0] _T_798 = _T_63 ? 2'h1 : _T_797; // @[Lookup.scala 33:37]
  wire [1:0] _T_799 = _T_61 ? 2'h1 : _T_798; // @[Lookup.scala 33:37]
  wire [1:0] _T_800 = _T_59 ? 2'h2 : _T_799; // @[Lookup.scala 33:37]
  wire [1:0] _T_801 = _T_57 ? 2'h2 : _T_800; // @[Lookup.scala 33:37]
  wire [1:0] _T_802 = _T_55 ? 2'h1 : _T_801; // @[Lookup.scala 33:37]
  wire [1:0] _T_803 = _T_53 ? 2'h1 : _T_802; // @[Lookup.scala 33:37]
  wire [1:0] _T_804 = _T_51 ? 2'h1 : _T_803; // @[Lookup.scala 33:37]
  wire [1:0] _T_805 = _T_49 ? 2'h1 : _T_804; // @[Lookup.scala 33:37]
  wire [1:0] _T_806 = _T_47 ? 2'h1 : _T_805; // @[Lookup.scala 33:37]
  wire [1:0] _T_807 = _T_45 ? 2'h1 : _T_806; // @[Lookup.scala 33:37]
  wire [1:0] _T_808 = _T_43 ? 2'h1 : _T_807; // @[Lookup.scala 33:37]
  wire [1:0] _T_809 = _T_41 ? 2'h1 : _T_808; // @[Lookup.scala 33:37]
  wire [1:0] _T_810 = _T_39 ? 2'h1 : _T_809; // @[Lookup.scala 33:37]
  wire [1:0] _T_811 = _T_37 ? 2'h1 : _T_810; // @[Lookup.scala 33:37]
  wire [1:0] csignals_5 = _T_35 ? 2'h2 : _T_811; // @[Lookup.scala 33:37]
  wire  _T_812 = ~csignals_0; // @[idu.scala 144:16]
  wire  _T_813 = fu_in_ex_et != 5'h0; // @[idu.scala 144:38]
  wire  has_ex = _T_812 | _T_813; // @[idu.scala 144:23]
  wire  _T_822 = ~io_ex_flush_valid; // @[idu.scala 159:37]
  wire [4:0] _T_827_et = _T_812 ? 5'h10 : 5'h0; // @[Mux.scala 87:16]
  wire [4:0] _T_827_code = _T_812 ? 5'ha : 5'h0; // @[Mux.scala 87:16]
  wire  _T_830 = ~_T_30; // @[idu.scala 176:31]
  wire  _T_831 = isu_io_fu_in_ready & isu_io_fu_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_832 = _T_830 & _T_831; // @[idu.scala 176:48]
  wire  _T_833 = io_ex_flush_valid | _T_832; // @[idu.scala 176:27]
  wire  _T_836 = _T_822 & _T_30; // @[idu.scala 178:34]
  wire  _GEN_6 = _T_836 | fu_valid; // @[idu.scala 178:54]
  ISU isu ( // @[idu.scala 21:19]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_fu_in_ready(isu_io_fu_in_ready),
    .io_fu_in_valid(isu_io_fu_in_valid),
    .io_fu_in_bits_pc(isu_io_fu_in_bits_pc),
    .io_fu_in_bits_instr_op(isu_io_fu_in_bits_instr_op),
    .io_fu_in_bits_instr_rs_idx(isu_io_fu_in_bits_instr_rs_idx),
    .io_fu_in_bits_instr_rt_idx(isu_io_fu_in_bits_instr_rt_idx),
    .io_fu_in_bits_instr_rd_idx(isu_io_fu_in_bits_instr_rd_idx),
    .io_fu_in_bits_instr_shamt(isu_io_fu_in_bits_instr_shamt),
    .io_fu_in_bits_instr_func(isu_io_fu_in_bits_instr_func),
    .io_fu_in_bits_fu_type(isu_io_fu_in_bits_fu_type),
    .io_fu_in_bits_fu_op(isu_io_fu_in_bits_fu_op),
    .io_fu_in_bits_op1_sel(isu_io_fu_in_bits_op1_sel),
    .io_fu_in_bits_op2_sel(isu_io_fu_in_bits_op2_sel),
    .io_fu_in_bits_opd_sel(isu_io_fu_in_bits_opd_sel),
    .io_fu_in_bits_ex_et(isu_io_fu_in_bits_ex_et),
    .io_fu_in_bits_ex_code(isu_io_fu_in_bits_ex_code),
    .io_fu_in_bits_ex_addr(isu_io_fu_in_bits_ex_addr),
    .io_fu_in_bits_ex_asid(isu_io_fu_in_bits_ex_asid),
    .io_fu_out_ready(isu_io_fu_out_ready),
    .io_fu_out_valid(isu_io_fu_out_valid),
    .io_fu_out_bits_wb_v(isu_io_fu_out_bits_wb_v),
    .io_fu_out_bits_wb_id(isu_io_fu_out_bits_wb_id),
    .io_fu_out_bits_wb_pc(isu_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(isu_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(isu_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(isu_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(isu_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(isu_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(isu_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_rd_idx(isu_io_fu_out_bits_wb_rd_idx),
    .io_fu_out_bits_wb_wen(isu_io_fu_out_bits_wb_wen),
    .io_fu_out_bits_wb_data(isu_io_fu_out_bits_wb_data),
    .io_fu_out_bits_wb_is_ds(isu_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_wb_is_br(isu_io_fu_out_bits_wb_is_br),
    .io_fu_out_bits_wb_npc(isu_io_fu_out_bits_wb_npc),
    .io_fu_out_bits_ops_fu_type(isu_io_fu_out_bits_ops_fu_type),
    .io_fu_out_bits_ops_fu_op(isu_io_fu_out_bits_ops_fu_op),
    .io_fu_out_bits_ops_op1(isu_io_fu_out_bits_ops_op1),
    .io_fu_out_bits_ops_op2(isu_io_fu_out_bits_ops_op2),
    .io_fu_out_bits_ex_et(isu_io_fu_out_bits_ex_et),
    .io_fu_out_bits_ex_code(isu_io_fu_out_bits_ex_code),
    .io_fu_out_bits_ex_addr(isu_io_fu_out_bits_ex_addr),
    .io_fu_out_bits_ex_asid(isu_io_fu_out_bits_ex_asid),
    .io_br_flush_valid(isu_io_br_flush_valid),
    .io_br_flush_bits_br_target(isu_io_br_flush_bits_br_target),
    .io_rfio_rs_idx(isu_io_rfio_rs_idx),
    .io_rfio_rt_idx(isu_io_rfio_rt_idx),
    .io_rfio_wen(isu_io_rfio_wen),
    .io_rfio_wid(isu_io_rfio_wid),
    .io_rfio_rd_idx(isu_io_rfio_rd_idx),
    .io_rfio_rs_data_valid(isu_io_rfio_rs_data_valid),
    .io_rfio_rs_data_bits(isu_io_rfio_rs_data_bits),
    .io_rfio_rt_data_valid(isu_io_rfio_rt_data_valid),
    .io_rfio_rt_data_bits(isu_io_rfio_rt_data_bits)
  );
  assign io_fu_in_ready = _T_32 | isu_io_fu_in_ready; // @[idu.scala 26:18]
  assign io_fu_out_valid = isu_io_fu_out_valid; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_v = isu_io_fu_out_bits_wb_v; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_id = isu_io_fu_out_bits_wb_id; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_pc = isu_io_fu_out_bits_wb_pc; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_instr_op = isu_io_fu_out_bits_wb_instr_op; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_instr_rs_idx = isu_io_fu_out_bits_wb_instr_rs_idx; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_instr_rt_idx = isu_io_fu_out_bits_wb_instr_rt_idx; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_instr_rd_idx = isu_io_fu_out_bits_wb_instr_rd_idx; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_instr_shamt = isu_io_fu_out_bits_wb_instr_shamt; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_instr_func = isu_io_fu_out_bits_wb_instr_func; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_rd_idx = isu_io_fu_out_bits_wb_rd_idx; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_wen = isu_io_fu_out_bits_wb_wen; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_data = isu_io_fu_out_bits_wb_data; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_is_ds = isu_io_fu_out_bits_wb_is_ds; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_is_br = isu_io_fu_out_bits_wb_is_br; // @[idu.scala 174:13]
  assign io_fu_out_bits_wb_npc = isu_io_fu_out_bits_wb_npc; // @[idu.scala 174:13]
  assign io_fu_out_bits_ops_fu_type = isu_io_fu_out_bits_ops_fu_type; // @[idu.scala 174:13]
  assign io_fu_out_bits_ops_fu_op = isu_io_fu_out_bits_ops_fu_op; // @[idu.scala 174:13]
  assign io_fu_out_bits_ops_op1 = isu_io_fu_out_bits_ops_op1; // @[idu.scala 174:13]
  assign io_fu_out_bits_ops_op2 = isu_io_fu_out_bits_ops_op2; // @[idu.scala 174:13]
  assign io_fu_out_bits_ex_et = isu_io_fu_out_bits_ex_et; // @[idu.scala 174:13]
  assign io_fu_out_bits_ex_code = isu_io_fu_out_bits_ex_code; // @[idu.scala 174:13]
  assign io_fu_out_bits_ex_addr = isu_io_fu_out_bits_ex_addr; // @[idu.scala 174:13]
  assign io_fu_out_bits_ex_asid = isu_io_fu_out_bits_ex_asid; // @[idu.scala 174:13]
  assign io_br_flush_valid = isu_io_br_flush_valid; // @[idu.scala 172:19]
  assign io_br_flush_bits_br_target = isu_io_br_flush_bits_br_target; // @[idu.scala 172:19]
  assign io_rfio_rs_idx = isu_io_rfio_rs_idx; // @[idu.scala 171:15]
  assign io_rfio_rt_idx = isu_io_rfio_rt_idx; // @[idu.scala 171:15]
  assign io_rfio_wen = isu_io_rfio_wen; // @[idu.scala 171:15]
  assign io_rfio_wid = isu_io_rfio_wid; // @[idu.scala 171:15]
  assign io_rfio_rd_idx = isu_io_rfio_rd_idx; // @[idu.scala 171:15]
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_fu_in_valid = fu_valid & _T_822; // @[idu.scala 159:22]
  assign isu_io_fu_in_bits_pc = fu_in_pc; // @[idu.scala 166:24]
  assign isu_io_fu_in_bits_instr_op = fu_in_instr[31:26]; // @[idu.scala 165:27]
  assign isu_io_fu_in_bits_instr_rs_idx = fu_in_instr[25:21]; // @[idu.scala 165:27]
  assign isu_io_fu_in_bits_instr_rt_idx = fu_in_instr[20:16]; // @[idu.scala 165:27]
  assign isu_io_fu_in_bits_instr_rd_idx = fu_in_instr[15:11]; // @[idu.scala 165:27]
  assign isu_io_fu_in_bits_instr_shamt = fu_in_instr[10:6]; // @[idu.scala 165:27]
  assign isu_io_fu_in_bits_instr_func = fu_in_instr[5:0]; // @[idu.scala 165:27]
  assign isu_io_fu_in_bits_fu_type = has_ex ? 3'h5 : csignals_1; // @[idu.scala 160:29]
  assign isu_io_fu_in_bits_fu_op = has_ex ? 5'h0 : csignals_2; // @[idu.scala 161:27]
  assign isu_io_fu_in_bits_op1_sel = has_ex ? 2'h0 : csignals_3; // @[idu.scala 162:29]
  assign isu_io_fu_in_bits_op2_sel = has_ex ? 3'h0 : csignals_4; // @[idu.scala 163:29]
  assign isu_io_fu_in_bits_opd_sel = has_ex ? 2'h0 : csignals_5; // @[idu.scala 164:29]
  assign isu_io_fu_in_bits_ex_et = _T_813 ? fu_in_ex_et : _T_827_et; // @[idu.scala 167:24]
  assign isu_io_fu_in_bits_ex_code = _T_813 ? fu_in_ex_code : _T_827_code; // @[idu.scala 167:24]
  assign isu_io_fu_in_bits_ex_addr = _T_813 ? fu_in_ex_addr : 32'h0; // @[idu.scala 167:24]
  assign isu_io_fu_in_bits_ex_asid = _T_813 ? fu_in_ex_asid : 8'h0; // @[idu.scala 167:24]
  assign isu_io_fu_out_ready = io_fu_out_ready; // @[idu.scala 174:13]
  assign isu_io_rfio_rs_data_valid = io_rfio_rs_data_valid; // @[idu.scala 171:15]
  assign isu_io_rfio_rs_data_bits = io_rfio_rs_data_bits; // @[idu.scala 171:15]
  assign isu_io_rfio_rt_data_valid = io_rfio_rt_data_valid; // @[idu.scala 171:15]
  assign isu_io_rfio_rt_data_bits = io_rfio_rt_data_bits; // @[idu.scala 171:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fu_in_pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fu_in_instr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  fu_in_ex_et = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fu_in_ex_code = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fu_in_ex_addr = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fu_in_ex_asid = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fu_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fu_in_pc <= 32'h0;
    end else if (_T_30) begin
      fu_in_pc <= io_fu_in_bits_pc;
    end
    if (reset) begin
      fu_in_instr <= 32'h0;
    end else if (_T_30) begin
      fu_in_instr <= io_fu_in_bits_instr;
    end
    if (reset) begin
      fu_in_ex_et <= 5'h0;
    end else if (_T_30) begin
      fu_in_ex_et <= io_fu_in_bits_ex_et;
    end
    if (reset) begin
      fu_in_ex_code <= 5'h0;
    end else if (_T_30) begin
      fu_in_ex_code <= io_fu_in_bits_ex_code;
    end
    if (reset) begin
      fu_in_ex_addr <= 32'h0;
    end else if (_T_30) begin
      fu_in_ex_addr <= io_fu_in_bits_ex_addr;
    end
    if (reset) begin
      fu_in_ex_asid <= 8'h0;
    end else if (_T_30) begin
      fu_in_ex_asid <= io_fu_in_bits_ex_asid;
    end
    if (reset) begin
      fu_valid <= 1'h0;
    end else if (_T_833) begin
      fu_valid <= 1'h0;
    end else begin
      fu_valid <= _GEN_6;
    end
  end
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input         io_fu_in_bits_wb_v,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_wen,
  input  [31:0] io_fu_in_bits_wb_data,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  input  [2:0]  io_fu_in_bits_ops_fu_type,
  input  [4:0]  io_fu_in_bits_ops_fu_op,
  input  [31:0] io_fu_in_bits_ops_op1,
  input  [31:0] io_fu_in_bits_ops_op2,
  input  [4:0]  io_fu_in_bits_ex_et,
  input  [4:0]  io_fu_in_bits_ex_code,
  input  [31:0] io_fu_in_bits_ex_addr,
  input  [7:0]  io_fu_in_bits_ex_asid,
  input         io_fu_out_ready,
  output        io_fu_out_valid,
  output        io_fu_out_bits_wb_v,
  output [7:0]  io_fu_out_bits_wb_id,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output [4:0]  io_fu_out_bits_wb_rd_idx,
  output        io_fu_out_bits_wb_wen,
  output [31:0] io_fu_out_bits_wb_data,
  output        io_fu_out_bits_wb_is_ds,
  output        io_fu_out_bits_wb_is_br,
  output [31:0] io_fu_out_bits_wb_npc,
  output [2:0]  io_fu_out_bits_ops_fu_type,
  output [4:0]  io_fu_out_bits_ops_fu_op,
  output [31:0] io_fu_out_bits_ops_op1,
  output [31:0] io_fu_out_bits_ops_op2,
  output [4:0]  io_fu_out_bits_ex_et,
  output [4:0]  io_fu_out_bits_ex_code,
  output [31:0] io_fu_out_bits_ex_addr,
  output [7:0]  io_fu_out_bits_ex_asid,
  output [31:0] io_cp0_rport_addr,
  input  [31:0] io_cp0_rport_data,
  output        io_cp0_wport_valid,
  output [31:0] io_cp0_wport_bits_addr,
  output [31:0] io_cp0_wport_bits_data,
  input  [4:0]  io_cp0_tlbr_port_index_index,
  input  [15:0] io_cp0_tlbr_port_pagemask_mask,
  input  [18:0] io_cp0_tlbr_port_entry_hi_vpn,
  input  [7:0]  io_cp0_tlbr_port_entry_hi_asid,
  input  [19:0] io_cp0_tlbr_port_entry_lo0_pfn,
  input  [2:0]  io_cp0_tlbr_port_entry_lo0_c,
  input         io_cp0_tlbr_port_entry_lo0_d,
  input         io_cp0_tlbr_port_entry_lo0_v,
  input         io_cp0_tlbr_port_entry_lo0_g,
  input  [19:0] io_cp0_tlbr_port_entry_lo1_pfn,
  input  [2:0]  io_cp0_tlbr_port_entry_lo1_c,
  input         io_cp0_tlbr_port_entry_lo1_d,
  input         io_cp0_tlbr_port_entry_lo1_v,
  input         io_cp0_tlbr_port_entry_lo1_g,
  output        io_cp0_tlbw_port_valid,
  output [15:0] io_cp0_tlbw_port_bits_pagemask_mask,
  output [18:0] io_cp0_tlbw_port_bits_entry_hi_vpn,
  output [7:0]  io_cp0_tlbw_port_bits_entry_hi_asid,
  output [19:0] io_cp0_tlbw_port_bits_entry_lo0_pfn,
  output [2:0]  io_cp0_tlbw_port_bits_entry_lo0_c,
  output        io_cp0_tlbw_port_bits_entry_lo0_d,
  output        io_cp0_tlbw_port_bits_entry_lo0_v,
  output        io_cp0_tlbw_port_bits_entry_lo0_g,
  output [19:0] io_cp0_tlbw_port_bits_entry_lo1_pfn,
  output [2:0]  io_cp0_tlbw_port_bits_entry_lo1_c,
  output        io_cp0_tlbw_port_bits_entry_lo1_d,
  output        io_cp0_tlbw_port_bits_entry_lo1_v,
  output        io_cp0_tlbw_port_bits_entry_lo1_g,
  output        io_cp0_tlbp_port_valid,
  output        io_cp0_tlbp_port_bits_index_p,
  output [4:0]  io_cp0_tlbp_port_bits_index_index,
  output        io_daddr_req_valid,
  output        io_daddr_req_bits_func,
  output [31:0] io_daddr_req_bits_vaddr,
  output [1:0]  io_daddr_req_bits_len,
  output        io_daddr_req_bits_is_aligned,
  input  [31:0] io_daddr_resp_bits_paddr,
  input  [4:0]  io_daddr_resp_bits_ex_et,
  input  [4:0]  io_daddr_resp_bits_ex_code,
  input  [31:0] io_daddr_resp_bits_ex_addr,
  input  [7:0]  io_daddr_resp_bits_ex_asid,
  output [4:0]  io_tlb_rport_index,
  input  [15:0] io_tlb_rport_entry_pagemask,
  input  [18:0] io_tlb_rport_entry_vpn,
  input         io_tlb_rport_entry_g,
  input  [7:0]  io_tlb_rport_entry_asid,
  input  [23:0] io_tlb_rport_entry_p0_pfn,
  input  [2:0]  io_tlb_rport_entry_p0_c,
  input         io_tlb_rport_entry_p0_d,
  input         io_tlb_rport_entry_p0_v,
  input  [23:0] io_tlb_rport_entry_p1_pfn,
  input  [2:0]  io_tlb_rport_entry_p1_c,
  input         io_tlb_rport_entry_p1_d,
  input         io_tlb_rport_entry_p1_v,
  output        io_tlb_wport_valid,
  output [4:0]  io_tlb_wport_bits_index,
  output [15:0] io_tlb_wport_bits_entry_pagemask,
  output [18:0] io_tlb_wport_bits_entry_vpn,
  output        io_tlb_wport_bits_entry_g,
  output [7:0]  io_tlb_wport_bits_entry_asid,
  output [23:0] io_tlb_wport_bits_entry_p0_pfn,
  output [2:0]  io_tlb_wport_bits_entry_p0_c,
  output        io_tlb_wport_bits_entry_p0_d,
  output        io_tlb_wport_bits_entry_p0_v,
  output [23:0] io_tlb_wport_bits_entry_p1_pfn,
  output [2:0]  io_tlb_wport_bits_entry_p1_c,
  output        io_tlb_wport_bits_entry_p1_d,
  output        io_tlb_wport_bits_entry_p1_v,
  output [18:0] io_tlb_pport_entry_hi_vpn,
  output [7:0]  io_tlb_pport_entry_hi_asid,
  input         io_tlb_pport_index_p,
  input  [4:0]  io_tlb_pport_index_index,
  output        io_icache_control_valid,
  output [2:0]  io_icache_control_bits_op,
  output [31:0] io_icache_control_bits_addr,
  output        io_bp_valid,
  output        io_bp_bits_v,
  output [4:0]  io_bp_bits_rd_idx,
  output        io_bp_bits_wen,
  output [31:0] io_bp_bits_data,
  input         io_ex_flush_valid
);
  wire  _T = io_fu_in_ready & io_fu_in_valid; // @[Decoupled.scala 40:37]
  reg  fu_in_wb_v; // @[Reg.scala 27:20]
  reg [31:0] _RAND_0;
  reg [7:0] fu_in_wb_id; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [31:0] fu_in_wb_pc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [5:0] fu_in_wb_instr_op; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [4:0] fu_in_wb_instr_rs_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [4:0] fu_in_wb_instr_rt_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [4:0] fu_in_wb_instr_rd_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [4:0] fu_in_wb_instr_shamt; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [5:0] fu_in_wb_instr_func; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [4:0] fu_in_wb_rd_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg  fu_in_wb_wen; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg [31:0] fu_in_wb_data; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg  fu_in_wb_is_ds; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg  fu_in_wb_is_br; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg [31:0] fu_in_wb_npc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg [2:0] fu_in_ops_fu_type; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg [4:0] fu_in_ops_fu_op; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg [31:0] fu_in_ops_op1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg [31:0] fu_in_ops_op2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  reg [4:0] fu_in_ex_et; // @[Reg.scala 27:20]
  reg [31:0] _RAND_19;
  reg [4:0] fu_in_ex_code; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  reg [31:0] fu_in_ex_addr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_21;
  reg [7:0] fu_in_ex_asid; // @[Reg.scala 27:20]
  reg [31:0] _RAND_22;
  reg  fu_valid; // @[exu.scala 36:25]
  reg [31:0] _RAND_23;
  wire  _T_2 = ~fu_valid; // @[exu.scala 38:41]
  wire  _T_3 = io_fu_out_ready | _T_2; // @[exu.scala 38:38]
  wire  _T_4 = ~io_ex_flush_valid; // @[exu.scala 38:55]
  wire [4:0] op2_sa = fu_in_ops_op2[4:0]; // @[exu.scala 44:20]
  wire  _T_6 = fu_in_ops_fu_op == 5'h0; // @[exu.scala 61:12]
  wire [31:0] _T_8 = fu_in_ops_op1 + fu_in_ops_op2; // @[exu.scala 61:34]
  wire  _T_9 = fu_in_ops_fu_op == 5'h1; // @[exu.scala 62:12]
  wire [31:0] _T_11 = fu_in_ops_op1 - fu_in_ops_op2; // @[exu.scala 62:34]
  wire  _T_12 = fu_in_ops_fu_op == 5'h2; // @[exu.scala 63:12]
  wire [62:0] _GEN_27 = {{31'd0}, fu_in_ops_op1}; // @[exu.scala 63:34]
  wire [62:0] _T_13 = _GEN_27 << op2_sa; // @[exu.scala 63:34]
  wire  _T_14 = fu_in_ops_fu_op == 5'h3; // @[exu.scala 64:12]
  wire [31:0] _T_15 = fu_in_ops_op1 >> op2_sa; // @[exu.scala 64:34]
  wire  _T_16 = fu_in_ops_fu_op == 5'h4; // @[exu.scala 65:12]
  wire [31:0] _T_19 = $signed(fu_in_ops_op1) >>> op2_sa; // @[exu.scala 65:52]
  wire  _T_20 = fu_in_ops_fu_op == 5'h5; // @[exu.scala 66:12]
  wire [31:0] _T_21 = fu_in_ops_op1 & fu_in_ops_op2; // @[exu.scala 66:34]
  wire  _T_22 = fu_in_ops_fu_op == 5'h6; // @[exu.scala 67:12]
  wire [31:0] _T_23 = fu_in_ops_op1 | fu_in_ops_op2; // @[exu.scala 67:34]
  wire  _T_24 = fu_in_ops_fu_op == 5'h7; // @[exu.scala 68:12]
  wire [31:0] _T_25 = fu_in_ops_op1 ^ fu_in_ops_op2; // @[exu.scala 68:34]
  wire  _T_26 = fu_in_ops_fu_op == 5'h8; // @[exu.scala 69:12]
  wire [31:0] _T_28 = ~_T_23; // @[exu.scala 69:29]
  wire  _T_29 = fu_in_ops_fu_op == 5'h9; // @[exu.scala 70:12]
  wire  _T_32 = $signed(fu_in_ops_op1) < $signed(fu_in_ops_op2); // @[exu.scala 70:41]
  wire  _T_33 = fu_in_ops_fu_op == 5'ha; // @[exu.scala 71:12]
  wire  _T_34 = fu_in_ops_op1 < fu_in_ops_op2; // @[exu.scala 71:34]
  wire  _T_35 = fu_in_ops_fu_op == 5'hb; // @[exu.scala 72:12]
  wire  _T_36 = fu_in_ops_fu_op == 5'hc; // @[exu.scala 73:12]
  wire  _T_37 = fu_in_ops_fu_op == 5'hd; // @[exu.scala 74:12]
  wire  _T_38 = fu_in_ops_fu_op == 5'he; // @[exu.scala 75:12]
  wire  _T_41 = fu_in_ops_fu_op == 5'hf; // @[exu.scala 76:12]
  wire  _T_44 = fu_in_ops_fu_op == 5'h10; // @[exu.scala 77:12]
  wire  _T_47 = fu_in_ops_op1[31:16] == 16'h0; // @[utils.scala 136:26]
  wire [15:0] _T_50 = _T_47 ? fu_in_ops_op1[15:0] : fu_in_ops_op1[31:16]; // @[utils.scala 138:20]
  wire  _T_52 = _T_50[15:8] == 8'h0; // @[utils.scala 139:28]
  wire [7:0] _T_55 = _T_52 ? _T_50[7:0] : _T_50[15:8]; // @[utils.scala 141:20]
  wire  _T_57 = _T_55[7:4] == 4'h0; // @[utils.scala 142:26]
  wire [3:0] _T_60 = _T_57 ? _T_55[3:0] : _T_55[7:4]; // @[utils.scala 144:20]
  wire  _T_62 = _T_60[3:2] == 2'h0; // @[utils.scala 145:26]
  wire  _T_64 = ~_T_60[1]; // @[utils.scala 147:27]
  wire  _T_66 = ~_T_60[3]; // @[utils.scala 147:37]
  wire  _T_67 = _T_62 ? _T_64 : _T_66; // @[utils.scala 147:18]
  wire  _T_68 = fu_in_ops_op1 == 32'h0; // @[utils.scala 149:12]
  wire [4:0] _T_72 = {_T_47,_T_52,_T_57,_T_62,_T_67}; // @[utils.scala 149:31]
  wire [5:0] _T_73 = _T_68 ? 6'h20 : {{1'd0}, _T_72}; // @[utils.scala 149:8]
  wire  _T_74 = fu_in_ops_fu_op == 5'h11; // @[exu.scala 78:12]
  wire  _T_78 = fu_in_ops_op1[31:16] == 16'hffff; // @[utils.scala 157:26]
  wire [15:0] _T_81 = _T_78 ? fu_in_ops_op1[15:0] : fu_in_ops_op1[31:16]; // @[utils.scala 159:20]
  wire  _T_84 = _T_81[15:8] == 8'hff; // @[utils.scala 160:28]
  wire [7:0] _T_87 = _T_84 ? _T_81[7:0] : _T_81[15:8]; // @[utils.scala 162:20]
  wire  _T_90 = _T_87[7:4] == 4'hf; // @[utils.scala 163:26]
  wire [3:0] _T_93 = _T_90 ? _T_87[3:0] : _T_87[7:4]; // @[utils.scala 165:20]
  wire  _T_96 = _T_93[3:2] == 2'h3; // @[utils.scala 166:26]
  wire  _T_99 = _T_96 ? _T_93[1] : _T_93[3]; // @[utils.scala 168:18]
  wire  _T_101 = fu_in_ops_op1 == 32'hffffffff; // @[utils.scala 170:12]
  wire [4:0] _T_105 = {_T_78,_T_84,_T_90,_T_96,_T_99}; // @[utils.scala 170:38]
  wire [5:0] _T_106 = _T_101 ? 6'h20 : {{1'd0}, _T_105}; // @[utils.scala 170:8]
  wire  _T_107 = fu_in_ops_fu_op == 5'h12; // @[exu.scala 79:12]
  wire [7:0] _T_110 = fu_in_ops_op1[7:0]; // @[exu.scala 79:47]
  wire [31:0] _T_111 = {{24{_T_110[7]}},_T_110}; // @[exu.scala 79:60]
  wire  _T_112 = fu_in_ops_fu_op == 5'h13; // @[exu.scala 80:12]
  wire [15:0] _T_115 = fu_in_ops_op1[15:0]; // @[exu.scala 80:48]
  wire [31:0] _T_116 = {{16{_T_115[15]}},_T_115}; // @[exu.scala 80:61]
  wire  _T_117 = fu_in_ops_fu_op == 5'h14; // @[exu.scala 81:12]
  wire [31:0] _T_124 = {fu_in_ops_op1[23:16],fu_in_ops_op1[31:24],fu_in_ops_op1[7:0],fu_in_ops_op1[15:8]}; // @[Cat.scala 29:58]
  wire  _T_125 = fu_in_ops_fu_op == 5'h15; // @[exu.scala 82:12]
  wire [4:0] _T_127 = fu_in_wb_instr_rd_idx - fu_in_wb_instr_shamt; // @[exu.scala 47:20]
  wire [5:0] _GEN_28 = {{1'd0}, _T_127}; // @[exu.scala 47:27]
  wire [5:0] _T_129 = _GEN_28 + 6'h1; // @[exu.scala 47:27]
  wire [63:0] _T_130 = 64'h1 << _T_129; // @[exu.scala 48:21]
  wire [63:0] _T_132 = _T_130 - 64'h1; // @[exu.scala 48:29]
  wire [94:0] _GEN_29 = {{31'd0}, _T_132}; // @[exu.scala 49:29]
  wire [94:0] _T_133 = _GEN_29 << fu_in_wb_instr_shamt; // @[exu.scala 49:29]
  wire [94:0] _T_134 = ~_T_133; // @[exu.scala 49:22]
  wire [94:0] _GEN_30 = {{63'd0}, fu_in_ops_op2}; // @[exu.scala 49:20]
  wire [94:0] _T_135 = _GEN_30 & _T_134; // @[exu.scala 49:20]
  wire [63:0] _GEN_31 = {{32'd0}, fu_in_ops_op1}; // @[exu.scala 49:46]
  wire [63:0] _T_136 = _GEN_31 & _T_132; // @[exu.scala 49:46]
  wire [94:0] _GEN_32 = {{31'd0}, _T_136}; // @[exu.scala 49:54]
  wire [94:0] _T_137 = _GEN_32 << fu_in_wb_instr_shamt; // @[exu.scala 49:54]
  wire [94:0] _T_138 = _T_135 | _T_137; // @[exu.scala 49:38]
  wire  _T_140 = fu_in_ops_fu_op == 5'h16; // @[exu.scala 83:12]
  wire [5:0] _GEN_33 = {{1'd0}, fu_in_wb_instr_rd_idx}; // @[exu.scala 54:20]
  wire [5:0] _T_142 = _GEN_33 + 6'h1; // @[exu.scala 54:20]
  wire [63:0] _T_143 = 64'h1 << _T_142; // @[exu.scala 55:21]
  wire [63:0] _T_145 = _T_143 - 64'h1; // @[exu.scala 55:30]
  wire [94:0] _GEN_34 = {{31'd0}, _T_145}; // @[exu.scala 56:29]
  wire [94:0] _T_146 = _GEN_34 << fu_in_wb_instr_shamt; // @[exu.scala 56:29]
  wire [94:0] _GEN_35 = {{63'd0}, fu_in_ops_op1}; // @[exu.scala 56:21]
  wire [94:0] _T_147 = _GEN_35 & _T_146; // @[exu.scala 56:21]
  wire [94:0] _T_148 = _T_147 >> fu_in_wb_instr_shamt; // @[exu.scala 56:38]
  wire  _T_150 = fu_in_ops_fu_op == 5'h17; // @[exu.scala 84:12]
  wire [5:0] _GEN_36 = {{1'd0}, op2_sa}; // @[exu.scala 84:62]
  wire [5:0] _T_153 = 6'h20 - _GEN_36; // @[exu.scala 84:62]
  wire [94:0] _T_154 = _GEN_35 << _T_153; // @[exu.scala 84:53]
  wire [94:0] _GEN_38 = {{63'd0}, _T_15}; // @[exu.scala 84:46]
  wire [94:0] _T_155 = _GEN_38 | _T_154; // @[exu.scala 84:46]
  wire [31:0] _T_156 = _T_6 ? _T_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_157 = _T_9 ? _T_11 : 32'h0; // @[Mux.scala 27:72]
  wire [62:0] _T_158 = _T_12 ? _T_13 : 63'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_159 = _T_14 ? _T_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_160 = _T_16 ? _T_19 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_161 = _T_20 ? _T_21 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_162 = _T_22 ? _T_23 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_163 = _T_24 ? _T_25 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_164 = _T_26 ? _T_28 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_165 = _T_29 & _T_32; // @[Mux.scala 27:72]
  wire  _T_166 = _T_33 & _T_34; // @[Mux.scala 27:72]
  wire [31:0] _T_167 = _T_35 ? fu_in_ops_op2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_168 = _T_36 ? fu_in_ops_op1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_169 = _T_37 ? fu_in_ops_op1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_170 = _T_38 ? _T_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_171 = _T_41 ? _T_11 : 32'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_172 = _T_44 ? _T_73 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_173 = _T_74 ? _T_106 : 6'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_174 = _T_107 ? _T_111 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_175 = _T_112 ? _T_116 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_176 = _T_117 ? _T_124 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_177 = _T_125 ? _T_138[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_178 = _T_140 ? _T_148[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [94:0] _T_179 = _T_150 ? _T_155 : 95'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_180 = _T_156 | _T_157; // @[Mux.scala 27:72]
  wire [62:0] _GEN_39 = {{31'd0}, _T_180}; // @[Mux.scala 27:72]
  wire [62:0] _T_181 = _GEN_39 | _T_158; // @[Mux.scala 27:72]
  wire [62:0] _GEN_40 = {{31'd0}, _T_159}; // @[Mux.scala 27:72]
  wire [62:0] _T_182 = _T_181 | _GEN_40; // @[Mux.scala 27:72]
  wire [62:0] _GEN_41 = {{31'd0}, _T_160}; // @[Mux.scala 27:72]
  wire [62:0] _T_183 = _T_182 | _GEN_41; // @[Mux.scala 27:72]
  wire [62:0] _GEN_42 = {{31'd0}, _T_161}; // @[Mux.scala 27:72]
  wire [62:0] _T_184 = _T_183 | _GEN_42; // @[Mux.scala 27:72]
  wire [62:0] _GEN_43 = {{31'd0}, _T_162}; // @[Mux.scala 27:72]
  wire [62:0] _T_185 = _T_184 | _GEN_43; // @[Mux.scala 27:72]
  wire [62:0] _GEN_44 = {{31'd0}, _T_163}; // @[Mux.scala 27:72]
  wire [62:0] _T_186 = _T_185 | _GEN_44; // @[Mux.scala 27:72]
  wire [62:0] _GEN_45 = {{31'd0}, _T_164}; // @[Mux.scala 27:72]
  wire [62:0] _T_187 = _T_186 | _GEN_45; // @[Mux.scala 27:72]
  wire [62:0] _GEN_46 = {{62'd0}, _T_165}; // @[Mux.scala 27:72]
  wire [62:0] _T_188 = _T_187 | _GEN_46; // @[Mux.scala 27:72]
  wire [62:0] _GEN_47 = {{62'd0}, _T_166}; // @[Mux.scala 27:72]
  wire [62:0] _T_189 = _T_188 | _GEN_47; // @[Mux.scala 27:72]
  wire [62:0] _GEN_48 = {{31'd0}, _T_167}; // @[Mux.scala 27:72]
  wire [62:0] _T_190 = _T_189 | _GEN_48; // @[Mux.scala 27:72]
  wire [62:0] _GEN_49 = {{31'd0}, _T_168}; // @[Mux.scala 27:72]
  wire [62:0] _T_191 = _T_190 | _GEN_49; // @[Mux.scala 27:72]
  wire [62:0] _GEN_50 = {{31'd0}, _T_169}; // @[Mux.scala 27:72]
  wire [62:0] _T_192 = _T_191 | _GEN_50; // @[Mux.scala 27:72]
  wire [62:0] _GEN_51 = {{31'd0}, _T_170}; // @[Mux.scala 27:72]
  wire [62:0] _T_193 = _T_192 | _GEN_51; // @[Mux.scala 27:72]
  wire [62:0] _GEN_52 = {{31'd0}, _T_171}; // @[Mux.scala 27:72]
  wire [62:0] _T_194 = _T_193 | _GEN_52; // @[Mux.scala 27:72]
  wire [62:0] _GEN_53 = {{57'd0}, _T_172}; // @[Mux.scala 27:72]
  wire [62:0] _T_195 = _T_194 | _GEN_53; // @[Mux.scala 27:72]
  wire [62:0] _GEN_54 = {{57'd0}, _T_173}; // @[Mux.scala 27:72]
  wire [62:0] _T_196 = _T_195 | _GEN_54; // @[Mux.scala 27:72]
  wire [62:0] _GEN_55 = {{31'd0}, _T_174}; // @[Mux.scala 27:72]
  wire [62:0] _T_197 = _T_196 | _GEN_55; // @[Mux.scala 27:72]
  wire [62:0] _GEN_56 = {{31'd0}, _T_175}; // @[Mux.scala 27:72]
  wire [62:0] _T_198 = _T_197 | _GEN_56; // @[Mux.scala 27:72]
  wire [62:0] _GEN_57 = {{31'd0}, _T_176}; // @[Mux.scala 27:72]
  wire [62:0] _T_199 = _T_198 | _GEN_57; // @[Mux.scala 27:72]
  wire [62:0] _GEN_58 = {{31'd0}, _T_177}; // @[Mux.scala 27:72]
  wire [62:0] _T_200 = _T_199 | _GEN_58; // @[Mux.scala 27:72]
  wire [62:0] _GEN_59 = {{31'd0}, _T_178}; // @[Mux.scala 27:72]
  wire [62:0] _T_201 = _T_200 | _GEN_59; // @[Mux.scala 27:72]
  wire [94:0] _GEN_60 = {{32'd0}, _T_201}; // @[Mux.scala 27:72]
  wire [94:0] _T_202 = _GEN_60 | _T_179; // @[Mux.scala 27:72]
  wire [31:0] alu_wdata = _T_202[31:0]; // @[exu.scala 85:5]
  wire  _T_206 = ~fu_in_ops_op1[31]; // @[exu.scala 87:34]
  wire  _T_208 = ~fu_in_ops_op2[31]; // @[exu.scala 87:46]
  wire  _T_209 = _T_206 & _T_208; // @[exu.scala 87:43]
  wire  _T_211 = _T_209 & alu_wdata[31]; // @[exu.scala 87:55]
  wire  _T_214 = fu_in_ops_op1[31] & fu_in_ops_op2[31]; // @[exu.scala 87:85]
  wire  _T_216 = ~alu_wdata[31]; // @[exu.scala 87:99]
  wire  _T_217 = _T_214 & _T_216; // @[exu.scala 87:96]
  wire  _T_218 = _T_211 | _T_217; // @[exu.scala 87:73]
  wire  _T_223 = _T_206 & fu_in_ops_op2[31]; // @[exu.scala 88:43]
  wire  _T_225 = _T_223 & alu_wdata[31]; // @[exu.scala 88:54]
  wire  _T_229 = fu_in_ops_op1[31] & _T_208; // @[exu.scala 88:84]
  wire  _T_232 = _T_229 & _T_216; // @[exu.scala 88:96]
  wire  _T_233 = _T_225 | _T_232; // @[exu.scala 88:72]
  wire  _T_234 = _T_38 & _T_218; // @[Mux.scala 27:72]
  wire  _T_235 = _T_41 & _T_233; // @[Mux.scala 27:72]
  wire  alu_ov = _T_234 | _T_235; // @[Mux.scala 27:72]
  wire  _T_237 = ~alu_ov; // @[exu.scala 89:25]
  wire  _T_239 = fu_in_ops_op2 != 32'h0; // @[exu.scala 90:34]
  wire  _T_241 = fu_in_ops_op2 == 32'h0; // @[exu.scala 91:34]
  wire  _T_242 = _T_37 ? _T_241 : _T_237; // @[Mux.scala 87:16]
  wire  alu_wen = _T_36 ? _T_239 : _T_242; // @[Mux.scala 87:16]
  wire [4:0] alu_ex_et = alu_ov ? 5'hc : 5'h0; // @[exu.scala 93:19]
  wire  _T_250 = io_fu_in_bits_ops_fu_type == 3'h3; // @[exu.scala 100:31]
  wire [7:0] cpr_addr = {fu_in_wb_instr_rd_idx,fu_in_wb_instr_func[2:0]}; // @[Cat.scala 29:58]
  wire  _T_253 = fu_in_ops_fu_type == 3'h5; // @[exu.scala 111:25]
  wire  pru_wen = _T_253 & _T_14; // @[exu.scala 111:36]
  wire  _T_255 = io_fu_out_ready & io_fu_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_257 = _T_255 & _T_253; // @[exu.scala 115:42]
  wire  _T_263 = $signed(fu_in_ops_op1) >= $signed(fu_in_ops_op2); // @[exu.scala 123:36]
  wire [1:0] _T_264 = {1'h1,_T_263}; // @[Cat.scala 29:58]
  wire  _T_265 = fu_in_ops_op1 >= fu_in_ops_op2; // @[exu.scala 124:29]
  wire [1:0] _T_266 = {1'h1,_T_265}; // @[Cat.scala 29:58]
  wire [1:0] _T_270 = {1'h1,_T_32}; // @[Cat.scala 29:58]
  wire [1:0] _T_272 = {1'h1,_T_34}; // @[Cat.scala 29:58]
  wire  _T_273 = fu_in_ops_op1 == fu_in_ops_op2; // @[exu.scala 127:29]
  wire [1:0] _T_274 = {1'h1,_T_273}; // @[Cat.scala 29:58]
  wire  _T_275 = fu_in_ops_op1 != fu_in_ops_op2; // @[exu.scala 128:29]
  wire [1:0] _T_276 = {1'h1,_T_275}; // @[Cat.scala 29:58]
  wire  _T_293 = 5'h18 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_294 = _T_293 ? _T_276 : 2'h0; // @[Mux.scala 68:16]
  wire  _T_295 = 5'h17 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_296 = _T_295 ? _T_274 : _T_294; // @[Mux.scala 68:16]
  wire  _T_297 = 5'h16 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_298 = _T_297 ? _T_272 : _T_296; // @[Mux.scala 68:16]
  wire  _T_299 = 5'h15 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_300 = _T_299 ? _T_270 : _T_298; // @[Mux.scala 68:16]
  wire  _T_301 = 5'h14 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_302 = _T_301 ? _T_266 : _T_300; // @[Mux.scala 68:16]
  wire  _T_303 = 5'h13 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_304 = _T_303 ? _T_264 : _T_302; // @[Mux.scala 68:16]
  wire  _T_305 = 5'h12 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_306 = _T_305 ? _T_276 : _T_304; // @[Mux.scala 68:16]
  wire  _T_307 = 5'h11 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_308 = _T_307 ? _T_274 : _T_306; // @[Mux.scala 68:16]
  wire  _T_309 = 5'h10 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_310 = _T_309 ? _T_272 : _T_308; // @[Mux.scala 68:16]
  wire  _T_311 = 5'hf == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_312 = _T_311 ? _T_270 : _T_310; // @[Mux.scala 68:16]
  wire  _T_313 = 5'he == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] _T_314 = _T_313 ? _T_266 : _T_312; // @[Mux.scala 68:16]
  wire  _T_315 = 5'hd == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [1:0] pru_trap = _T_315 ? _T_264 : _T_314; // @[Mux.scala 68:16]
  wire  _T_316 = 5'h2 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [4:0] _T_317 = _T_316 ? 5'h16 : fu_in_ex_et; // @[Mux.scala 68:16]
  wire  _T_318 = 5'h9 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [4:0] _T_319 = _T_318 ? 5'hf : _T_317; // @[Mux.scala 68:16]
  wire  _T_320 = 5'h1 == fu_in_ops_fu_op; // @[Mux.scala 68:19]
  wire [4:0] pru_normal_et = _T_320 ? 5'he : _T_319; // @[Mux.scala 68:16]
  wire [4:0] _T_322 = _T_318 ? 5'h9 : fu_in_ex_code; // @[Mux.scala 68:16]
  wire [4:0] pru_normal_code = _T_320 ? 5'h8 : _T_322; // @[Mux.scala 68:16]
  wire [4:0] _T_326 = pru_trap[0] ? 5'hd : 5'h0; // @[exu.scala 144:36]
  wire [4:0] pru_ex_et = pru_trap[1] ? _T_326 : pru_normal_et; // @[exu.scala 144:19]
  wire [4:0] pru_ex_code = pru_trap[1] ? _T_326 : pru_normal_code; // @[exu.scala 146:21]
  wire  _T_332 = 3'h5 == fu_in_ops_fu_type; // @[Mux.scala 68:19]
  wire [4:0] _T_333_et = _T_332 ? pru_ex_et : fu_in_ex_et; // @[Mux.scala 68:16]
  wire [4:0] _T_333_code = _T_332 ? pru_ex_code : fu_in_ex_code; // @[Mux.scala 68:16]
  wire  _T_334 = 3'h3 == fu_in_ops_fu_type; // @[Mux.scala 68:19]
  wire [4:0] _T_335_et = _T_334 ? io_daddr_resp_bits_ex_et : _T_333_et; // @[Mux.scala 68:16]
  wire [4:0] _T_335_code = _T_334 ? io_daddr_resp_bits_ex_code : _T_333_code; // @[Mux.scala 68:16]
  wire [31:0] _T_335_addr = _T_334 ? io_daddr_resp_bits_ex_addr : fu_in_ex_addr; // @[Mux.scala 68:16]
  wire [7:0] _T_335_asid = _T_334 ? io_daddr_resp_bits_ex_asid : fu_in_ex_asid; // @[Mux.scala 68:16]
  wire  _T_336 = 3'h1 == fu_in_ops_fu_type; // @[Mux.scala 68:19]
  wire [33:0] _T_339 = {fu_in_wb_v,fu_in_wb_wen,fu_in_wb_data}; // @[Cat.scala 29:58]
  wire [33:0] _T_341 = {1'h1,alu_wen,alu_wdata}; // @[Cat.scala 29:58]
  wire [33:0] _T_343 = {pru_wen,pru_wen,io_cp0_rport_data}; // @[Cat.scala 29:58]
  wire [33:0] _T_345 = _T_332 ? _T_343 : _T_339; // @[Mux.scala 68:16]
  wire [33:0] wb_info = _T_336 ? _T_341 : _T_345; // @[Mux.scala 68:16]
  wire  _T_350 = fu_in_ops_fu_type == 3'h3; // @[exu.scala 164:51]
  wire  _T_353 = io_daddr_resp_bits_ex_et != 5'h0; // @[exu.scala 167:15]
  wire [2:0] _T_354 = _T_353 ? 3'h5 : 3'h3; // @[exu.scala 166:70]
  wire [1:0] cache_control_target = fu_in_ops_op2[1:0]; // @[exu.scala 178:43]
  wire  _T_360 = _T_257 & _T_33; // @[exu.scala 181:24]
  wire  _T_361 = cache_control_target == 2'h0; // @[exu.scala 182:26]
  wire [31:0] tlbr_mask = {{16'd0}, io_tlb_rport_entry_pagemask}; // @[exu.scala 187:55 exu.scala 187:55]
  wire [31:0] _T_368 = ~tlbr_mask; // @[exu.scala 194:66]
  wire [31:0] _GEN_61 = {{13'd0}, io_tlb_rport_entry_vpn}; // @[exu.scala 194:64]
  wire [31:0] _T_369 = _GEN_61 & _T_368; // @[exu.scala 194:64]
  wire [31:0] _GEN_62 = {{24'd0}, io_tlb_rport_entry_asid}; // @[exu.scala 195:66]
  wire [31:0] _T_371 = _GEN_62 & _T_368; // @[exu.scala 195:66]
  wire [31:0] _GEN_63 = {{8'd0}, io_tlb_rport_entry_p0_pfn}; // @[exu.scala 201:68]
  wire [31:0] _T_373 = _GEN_63 & _T_368; // @[exu.scala 201:68]
  wire [31:0] _GEN_64 = {{8'd0}, io_tlb_rport_entry_p1_pfn}; // @[exu.scala 208:68]
  wire [31:0] _T_375 = _GEN_64 & _T_368; // @[exu.scala 208:68]
  reg [4:0] cpr_random_index; // @[exu.scala 213:27]
  reg [31:0] _RAND_24;
  wire [31:0] _T_377 = {{16'd0}, io_cp0_tlbr_port_pagemask_mask}; // @[exu.scala 214:59 exu.scala 214:59]
  wire [31:0] tlbw_mask = ~_T_377; // @[exu.scala 214:19]
  wire  _T_383 = _T_22 | _T_24; // @[exu.scala 216:48]
  wire [31:0] _GEN_65 = {{13'd0}, io_cp0_tlbr_port_entry_hi_vpn}; // @[exu.scala 220:64]
  wire [31:0] _T_387 = _GEN_65 & tlbw_mask; // @[exu.scala 220:64]
  wire [31:0] _GEN_66 = {{12'd0}, io_cp0_tlbr_port_entry_lo0_pfn}; // @[exu.scala 223:68]
  wire [31:0] _T_389 = _GEN_66 & tlbw_mask; // @[exu.scala 223:68]
  wire [31:0] _GEN_67 = {{12'd0}, io_cp0_tlbr_port_entry_lo1_pfn}; // @[exu.scala 227:68]
  wire [31:0] _T_390 = _GEN_67 & tlbw_mask; // @[exu.scala 227:68]
  wire  _T_392 = io_tlb_wport_valid & _T_24; // @[exu.scala 231:28]
  wire  _T_394 = _T_392 & _T_4; // @[exu.scala 231:51]
  wire [4:0] _T_396 = cpr_random_index + 5'h1; // @[exu.scala 232:42]
  wire  _T_403 = ~_T; // @[exu.scala 242:31]
  wire  _T_405 = _T_403 & _T_255; // @[exu.scala 242:48]
  wire  _T_406 = io_ex_flush_valid | _T_405; // @[exu.scala 242:27]
  wire  _T_409 = _T_4 & _T; // @[exu.scala 244:34]
  wire  _GEN_25 = _T_409 | fu_valid; // @[exu.scala 244:54]
  assign io_fu_in_ready = _T_3 & _T_4; // @[exu.scala 38:18]
  assign io_fu_out_valid = fu_valid; // @[exu.scala 154:19]
  assign io_fu_out_bits_wb_v = wb_info[33]; // @[exu.scala 155:21 exu.scala 160:23]
  assign io_fu_out_bits_wb_id = fu_in_wb_id; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_pc = fu_in_wb_pc; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_instr_op = fu_in_wb_instr_op; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_instr_rs_idx = fu_in_wb_instr_rs_idx; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_instr_rt_idx = fu_in_wb_instr_rt_idx; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_instr_rd_idx = fu_in_wb_instr_rd_idx; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_instr_shamt = fu_in_wb_instr_shamt; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_instr_func = fu_in_wb_instr_func; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_rd_idx = fu_in_wb_rd_idx; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_wen = wb_info[32]; // @[exu.scala 155:21 exu.scala 161:25]
  assign io_fu_out_bits_wb_data = wb_info[31:0]; // @[exu.scala 155:21 exu.scala 162:26]
  assign io_fu_out_bits_wb_is_ds = fu_in_wb_is_ds; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_is_br = fu_in_wb_is_br; // @[exu.scala 155:21]
  assign io_fu_out_bits_wb_npc = fu_in_wb_npc; // @[exu.scala 155:21]
  assign io_fu_out_bits_ops_fu_type = _T_350 ? _T_354 : fu_in_ops_fu_type; // @[exu.scala 163:22 exu.scala 166:30]
  assign io_fu_out_bits_ops_fu_op = fu_in_ops_fu_op; // @[exu.scala 163:22]
  assign io_fu_out_bits_ops_op1 = _T_350 ? io_daddr_resp_bits_paddr : fu_in_ops_op1; // @[exu.scala 163:22 exu.scala 164:26]
  assign io_fu_out_bits_ops_op2 = fu_in_ops_op2; // @[exu.scala 163:22]
  assign io_fu_out_bits_ex_et = _T_336 ? alu_ex_et : _T_335_et; // @[exu.scala 150:21]
  assign io_fu_out_bits_ex_code = _T_336 ? 5'hc : _T_335_code; // @[exu.scala 150:21]
  assign io_fu_out_bits_ex_addr = _T_336 ? 32'h0 : _T_335_addr; // @[exu.scala 150:21]
  assign io_fu_out_bits_ex_asid = _T_336 ? 8'h0 : _T_335_asid; // @[exu.scala 150:21]
  assign io_cp0_rport_addr = {{24'd0}, cpr_addr}; // @[exu.scala 110:21]
  assign io_cp0_wport_valid = _T_257 & _T_16; // @[exu.scala 115:22]
  assign io_cp0_wport_bits_addr = {{24'd0}, cpr_addr}; // @[exu.scala 117:26]
  assign io_cp0_wport_bits_data = fu_in_ops_op1; // @[exu.scala 118:26]
  assign io_cp0_tlbw_port_valid = _T_257 & _T_20; // @[exu.scala 189:26]
  assign io_cp0_tlbw_port_bits_pagemask_mask = tlbr_mask[15:0]; // @[exu.scala 193:39]
  assign io_cp0_tlbw_port_bits_entry_hi_vpn = _T_369[18:0]; // @[exu.scala 194:38]
  assign io_cp0_tlbw_port_bits_entry_hi_asid = _T_371[7:0]; // @[exu.scala 195:39]
  assign io_cp0_tlbw_port_bits_entry_lo0_pfn = _T_373[19:0]; // @[exu.scala 201:39]
  assign io_cp0_tlbw_port_bits_entry_lo0_c = io_tlb_rport_entry_p0_c; // @[exu.scala 198:37]
  assign io_cp0_tlbw_port_bits_entry_lo0_d = io_tlb_rport_entry_p0_d; // @[exu.scala 199:37]
  assign io_cp0_tlbw_port_bits_entry_lo0_v = io_tlb_rport_entry_p0_v; // @[exu.scala 197:37]
  assign io_cp0_tlbw_port_bits_entry_lo0_g = io_tlb_rport_entry_g; // @[exu.scala 200:37]
  assign io_cp0_tlbw_port_bits_entry_lo1_pfn = _T_375[19:0]; // @[exu.scala 208:39]
  assign io_cp0_tlbw_port_bits_entry_lo1_c = io_tlb_rport_entry_p1_c; // @[exu.scala 205:37]
  assign io_cp0_tlbw_port_bits_entry_lo1_d = io_tlb_rport_entry_p1_d; // @[exu.scala 206:37]
  assign io_cp0_tlbw_port_bits_entry_lo1_v = io_tlb_rport_entry_p1_v; // @[exu.scala 204:37]
  assign io_cp0_tlbw_port_bits_entry_lo1_g = io_tlb_rport_entry_g; // @[exu.scala 207:37]
  assign io_cp0_tlbp_port_valid = _T_257 & _T_26; // @[exu.scala 237:26]
  assign io_cp0_tlbp_port_bits_index_p = io_tlb_pport_index_p; // @[exu.scala 239:31]
  assign io_cp0_tlbp_port_bits_index_index = io_tlb_pport_index_index; // @[exu.scala 239:31]
  assign io_daddr_req_valid = _T & _T_250; // @[exu.scala 99:22]
  assign io_daddr_req_bits_func = io_fu_in_bits_ops_fu_op[3]; // @[exu.scala 102:26]
  assign io_daddr_req_bits_vaddr = io_fu_in_bits_ops_op1; // @[exu.scala 101:27]
  assign io_daddr_req_bits_len = io_fu_in_bits_ops_fu_op[2:1]; // @[exu.scala 103:25]
  assign io_daddr_req_bits_is_aligned = io_fu_in_bits_ops_fu_op[4]; // @[exu.scala 104:32]
  assign io_tlb_rport_index = io_cp0_tlbr_port_index_index; // @[exu.scala 188:22]
  assign io_tlb_wport_valid = _T_257 & _T_383; // @[exu.scala 215:22]
  assign io_tlb_wport_bits_index = _T_22 ? io_cp0_tlbr_port_index_index : cpr_random_index; // @[exu.scala 218:27]
  assign io_tlb_wport_bits_entry_pagemask = io_cp0_tlbr_port_pagemask_mask; // @[exu.scala 219:36]
  assign io_tlb_wport_bits_entry_vpn = _T_387[18:0]; // @[exu.scala 220:31]
  assign io_tlb_wport_bits_entry_g = io_cp0_tlbr_port_entry_lo0_g & io_cp0_tlbr_port_entry_lo1_g; // @[exu.scala 222:29]
  assign io_tlb_wport_bits_entry_asid = io_cp0_tlbr_port_entry_hi_asid; // @[exu.scala 221:32]
  assign io_tlb_wport_bits_entry_p0_pfn = _T_389[23:0]; // @[exu.scala 223:34]
  assign io_tlb_wport_bits_entry_p0_c = io_cp0_tlbr_port_entry_lo0_c; // @[exu.scala 224:32]
  assign io_tlb_wport_bits_entry_p0_d = io_cp0_tlbr_port_entry_lo0_d; // @[exu.scala 225:32]
  assign io_tlb_wport_bits_entry_p0_v = io_cp0_tlbr_port_entry_lo0_v; // @[exu.scala 226:32]
  assign io_tlb_wport_bits_entry_p1_pfn = _T_390[23:0]; // @[exu.scala 227:34]
  assign io_tlb_wport_bits_entry_p1_c = io_cp0_tlbr_port_entry_lo1_c; // @[exu.scala 228:32]
  assign io_tlb_wport_bits_entry_p1_d = io_cp0_tlbr_port_entry_lo1_d; // @[exu.scala 229:32]
  assign io_tlb_wport_bits_entry_p1_v = io_cp0_tlbr_port_entry_lo1_v; // @[exu.scala 230:32]
  assign io_tlb_pport_entry_hi_vpn = io_cp0_tlbr_port_entry_hi_vpn; // @[exu.scala 236:25]
  assign io_tlb_pport_entry_hi_asid = io_cp0_tlbr_port_entry_hi_asid; // @[exu.scala 236:25]
  assign io_icache_control_valid = _T_360 & _T_361; // @[exu.scala 180:27]
  assign io_icache_control_bits_op = fu_in_ops_op2[4:2]; // @[exu.scala 183:29]
  assign io_icache_control_bits_addr = fu_in_ops_op1; // @[exu.scala 184:31]
  assign io_bp_valid = io_fu_out_valid; // @[exu.scala 171:15]
  assign io_bp_bits_v = io_fu_out_bits_wb_v; // @[exu.scala 172:16]
  assign io_bp_bits_rd_idx = io_fu_out_bits_wb_rd_idx; // @[exu.scala 173:21]
  assign io_bp_bits_wen = io_fu_out_bits_wb_wen; // @[exu.scala 174:18]
  assign io_bp_bits_data = io_fu_out_bits_wb_data; // @[exu.scala 175:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fu_in_wb_v = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fu_in_wb_id = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  fu_in_wb_pc = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fu_in_wb_instr_op = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fu_in_wb_instr_rs_idx = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fu_in_wb_instr_rt_idx = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fu_in_wb_instr_rd_idx = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  fu_in_wb_instr_shamt = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fu_in_wb_instr_func = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fu_in_wb_rd_idx = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fu_in_wb_wen = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fu_in_wb_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fu_in_wb_is_ds = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fu_in_wb_is_br = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fu_in_wb_npc = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fu_in_ops_fu_type = _RAND_15[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  fu_in_ops_fu_op = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  fu_in_ops_op1 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  fu_in_ops_op2 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  fu_in_ex_et = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  fu_in_ex_code = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  fu_in_ex_addr = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  fu_in_ex_asid = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  fu_valid = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  cpr_random_index = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fu_in_wb_v <= 1'h0;
    end else if (_T) begin
      fu_in_wb_v <= io_fu_in_bits_wb_v;
    end
    if (reset) begin
      fu_in_wb_id <= 8'h0;
    end else if (_T) begin
      fu_in_wb_id <= io_fu_in_bits_wb_id;
    end
    if (reset) begin
      fu_in_wb_pc <= 32'h0;
    end else if (_T) begin
      fu_in_wb_pc <= io_fu_in_bits_wb_pc;
    end
    if (reset) begin
      fu_in_wb_instr_op <= 6'h0;
    end else if (_T) begin
      fu_in_wb_instr_op <= io_fu_in_bits_wb_instr_op;
    end
    if (reset) begin
      fu_in_wb_instr_rs_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rs_idx <= io_fu_in_bits_wb_instr_rs_idx;
    end
    if (reset) begin
      fu_in_wb_instr_rt_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rt_idx <= io_fu_in_bits_wb_instr_rt_idx;
    end
    if (reset) begin
      fu_in_wb_instr_rd_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rd_idx <= io_fu_in_bits_wb_instr_rd_idx;
    end
    if (reset) begin
      fu_in_wb_instr_shamt <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_shamt <= io_fu_in_bits_wb_instr_shamt;
    end
    if (reset) begin
      fu_in_wb_instr_func <= 6'h0;
    end else if (_T) begin
      fu_in_wb_instr_func <= io_fu_in_bits_wb_instr_func;
    end
    if (reset) begin
      fu_in_wb_rd_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_rd_idx <= io_fu_in_bits_wb_rd_idx;
    end
    if (reset) begin
      fu_in_wb_wen <= 1'h0;
    end else if (_T) begin
      fu_in_wb_wen <= io_fu_in_bits_wb_wen;
    end
    if (reset) begin
      fu_in_wb_data <= 32'h0;
    end else if (_T) begin
      fu_in_wb_data <= io_fu_in_bits_wb_data;
    end
    if (reset) begin
      fu_in_wb_is_ds <= 1'h0;
    end else if (_T) begin
      fu_in_wb_is_ds <= io_fu_in_bits_wb_is_ds;
    end
    if (reset) begin
      fu_in_wb_is_br <= 1'h0;
    end else if (_T) begin
      fu_in_wb_is_br <= io_fu_in_bits_wb_is_br;
    end
    if (reset) begin
      fu_in_wb_npc <= 32'h0;
    end else if (_T) begin
      fu_in_wb_npc <= io_fu_in_bits_wb_npc;
    end
    if (reset) begin
      fu_in_ops_fu_type <= 3'h0;
    end else if (_T) begin
      fu_in_ops_fu_type <= io_fu_in_bits_ops_fu_type;
    end
    if (reset) begin
      fu_in_ops_fu_op <= 5'h0;
    end else if (_T) begin
      fu_in_ops_fu_op <= io_fu_in_bits_ops_fu_op;
    end
    if (reset) begin
      fu_in_ops_op1 <= 32'h0;
    end else if (_T) begin
      fu_in_ops_op1 <= io_fu_in_bits_ops_op1;
    end
    if (reset) begin
      fu_in_ops_op2 <= 32'h0;
    end else if (_T) begin
      fu_in_ops_op2 <= io_fu_in_bits_ops_op2;
    end
    if (reset) begin
      fu_in_ex_et <= 5'h0;
    end else if (_T) begin
      fu_in_ex_et <= io_fu_in_bits_ex_et;
    end
    if (reset) begin
      fu_in_ex_code <= 5'h0;
    end else if (_T) begin
      fu_in_ex_code <= io_fu_in_bits_ex_code;
    end
    if (reset) begin
      fu_in_ex_addr <= 32'h0;
    end else if (_T) begin
      fu_in_ex_addr <= io_fu_in_bits_ex_addr;
    end
    if (reset) begin
      fu_in_ex_asid <= 8'h0;
    end else if (_T) begin
      fu_in_ex_asid <= io_fu_in_bits_ex_asid;
    end
    if (reset) begin
      fu_valid <= 1'h0;
    end else if (_T_406) begin
      fu_valid <= 1'h0;
    end else begin
      fu_valid <= _GEN_25;
    end
    if (reset) begin
      cpr_random_index <= 5'h0;
    end else if (_T_394) begin
      cpr_random_index <= _T_396;
    end
  end
endmodule
module EHU(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input         io_fu_in_bits_wb_v,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_wen,
  input  [31:0] io_fu_in_bits_wb_data,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  input  [2:0]  io_fu_in_bits_ops_fu_type,
  input  [4:0]  io_fu_in_bits_ops_fu_op,
  input  [31:0] io_fu_in_bits_ops_op1,
  input  [31:0] io_fu_in_bits_ops_op2,
  input  [4:0]  io_fu_in_bits_ex_et,
  input  [4:0]  io_fu_in_bits_ex_code,
  input  [31:0] io_fu_in_bits_ex_addr,
  input  [7:0]  io_fu_in_bits_ex_asid,
  input         io_fu_out_ready,
  output        io_fu_out_valid,
  output        io_fu_out_bits_wb_v,
  output [7:0]  io_fu_out_bits_wb_id,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output [4:0]  io_fu_out_bits_wb_rd_idx,
  output        io_fu_out_bits_wb_wen,
  output [31:0] io_fu_out_bits_wb_data,
  output        io_fu_out_bits_wb_ip7,
  output        io_fu_out_bits_wb_is_ds,
  output        io_fu_out_bits_wb_is_br,
  output [31:0] io_fu_out_bits_wb_npc,
  output [2:0]  io_fu_out_bits_ops_fu_type,
  output [4:0]  io_fu_out_bits_ops_fu_op,
  output [31:0] io_fu_out_bits_ops_op1,
  output [31:0] io_fu_out_bits_ops_op2,
  output        io_fu_out_bits_is_cached,
  output        io_cp0_valid,
  input         io_cp0_ip7,
  output [4:0]  io_cp0_ex_et,
  output [4:0]  io_cp0_ex_code,
  output [31:0] io_cp0_ex_addr,
  output [7:0]  io_cp0_ex_asid,
  output [31:0] io_cp0_wb_pc,
  output        io_cp0_wb_is_ds,
  output        io_cp0_wb_is_br,
  output [31:0] io_cp0_wb_npc,
  input         io_ex_flush_valid
);
  reg  fu_valid; // @[ehu.scala 20:25]
  reg [31:0] _RAND_0;
  wire  _T = io_fu_in_ready & io_fu_in_valid; // @[Decoupled.scala 40:37]
  reg  fu_in_wb_v; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [7:0] fu_in_wb_id; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [31:0] fu_in_wb_pc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [5:0] fu_in_wb_instr_op; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [4:0] fu_in_wb_instr_rs_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [4:0] fu_in_wb_instr_rt_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [4:0] fu_in_wb_instr_rd_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [4:0] fu_in_wb_instr_shamt; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [5:0] fu_in_wb_instr_func; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg [4:0] fu_in_wb_rd_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg  fu_in_wb_wen; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg [31:0] fu_in_wb_data; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg  fu_in_wb_is_ds; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg  fu_in_wb_is_br; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg [31:0] fu_in_wb_npc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg [2:0] fu_in_ops_fu_type; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg [4:0] fu_in_ops_fu_op; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg [31:0] fu_in_ops_op1; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  reg [31:0] fu_in_ops_op2; // @[Reg.scala 27:20]
  reg [31:0] _RAND_19;
  reg  fu_in_is_cached; // @[Reg.scala 27:20]
  reg [31:0] _RAND_20;
  reg [4:0] fu_in_ex_et; // @[Reg.scala 27:20]
  reg [31:0] _RAND_21;
  reg [4:0] fu_in_ex_code; // @[Reg.scala 27:20]
  reg [31:0] _RAND_22;
  reg [31:0] fu_in_ex_addr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_23;
  reg [7:0] fu_in_ex_asid; // @[Reg.scala 27:20]
  reg [31:0] _RAND_24;
  wire  _GEN_4 = _T | fu_in_is_cached; // @[Reg.scala 28:19]
  wire  _T_2 = ~fu_valid; // @[ehu.scala 22:22]
  wire  _T_3 = _T_2 | io_fu_out_ready; // @[ehu.scala 22:32]
  wire  _T_4 = ~io_ex_flush_valid; // @[ehu.scala 22:55]
  wire  _T_6 = io_fu_out_ready & io_fu_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = ~_T; // @[ehu.scala 35:9]
  wire  _T_10 = _T_8 & _T_6; // @[ehu.scala 35:26]
  wire  _GEN_25 = _T | fu_valid; // @[ehu.scala 37:33]
  assign io_fu_in_ready = _T_3 & _T_4; // @[ehu.scala 22:18]
  assign io_fu_out_valid = fu_valid; // @[ehu.scala 24:19]
  assign io_fu_out_bits_wb_v = fu_in_wb_v; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_id = fu_in_wb_id; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_pc = fu_in_wb_pc; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_instr_op = fu_in_wb_instr_op; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_instr_rs_idx = fu_in_wb_instr_rs_idx; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_instr_rt_idx = fu_in_wb_instr_rt_idx; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_instr_rd_idx = fu_in_wb_instr_rd_idx; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_instr_shamt = fu_in_wb_instr_shamt; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_instr_func = fu_in_wb_instr_func; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_rd_idx = fu_in_wb_rd_idx; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_wen = fu_in_wb_wen; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_data = fu_in_wb_data; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_ip7 = io_cp0_ip7; // @[ehu.scala 25:21 ehu.scala 28:25]
  assign io_fu_out_bits_wb_is_ds = fu_in_wb_is_ds; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_is_br = fu_in_wb_is_br; // @[ehu.scala 25:21]
  assign io_fu_out_bits_wb_npc = fu_in_wb_npc; // @[ehu.scala 25:21]
  assign io_fu_out_bits_ops_fu_type = fu_in_ops_fu_type; // @[ehu.scala 26:22]
  assign io_fu_out_bits_ops_fu_op = fu_in_ops_fu_op; // @[ehu.scala 26:22]
  assign io_fu_out_bits_ops_op1 = fu_in_ops_op1; // @[ehu.scala 26:22]
  assign io_fu_out_bits_ops_op2 = fu_in_ops_op2; // @[ehu.scala 26:22]
  assign io_fu_out_bits_is_cached = fu_in_is_cached; // @[ehu.scala 27:28]
  assign io_cp0_valid = io_fu_out_ready & io_fu_out_valid; // @[ehu.scala 31:16]
  assign io_cp0_ex_et = fu_in_ex_et; // @[ehu.scala 33:13]
  assign io_cp0_ex_code = fu_in_ex_code; // @[ehu.scala 33:13]
  assign io_cp0_ex_addr = fu_in_ex_addr; // @[ehu.scala 33:13]
  assign io_cp0_ex_asid = fu_in_ex_asid; // @[ehu.scala 33:13]
  assign io_cp0_wb_pc = io_fu_out_bits_wb_pc; // @[ehu.scala 32:13]
  assign io_cp0_wb_is_ds = io_fu_out_bits_wb_is_ds; // @[ehu.scala 32:13]
  assign io_cp0_wb_is_br = io_fu_out_bits_wb_is_br; // @[ehu.scala 32:13]
  assign io_cp0_wb_npc = io_fu_out_bits_wb_npc; // @[ehu.scala 32:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fu_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fu_in_wb_v = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  fu_in_wb_id = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fu_in_wb_pc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fu_in_wb_instr_op = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fu_in_wb_instr_rs_idx = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fu_in_wb_instr_rt_idx = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  fu_in_wb_instr_rd_idx = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fu_in_wb_instr_shamt = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fu_in_wb_instr_func = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fu_in_wb_rd_idx = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fu_in_wb_wen = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fu_in_wb_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fu_in_wb_is_ds = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fu_in_wb_is_br = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fu_in_wb_npc = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  fu_in_ops_fu_type = _RAND_16[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  fu_in_ops_fu_op = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  fu_in_ops_op1 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  fu_in_ops_op2 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  fu_in_is_cached = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  fu_in_ex_et = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  fu_in_ex_code = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  fu_in_ex_addr = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  fu_in_ex_asid = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fu_valid <= 1'h0;
    end else if (_T_10) begin
      fu_valid <= 1'h0;
    end else begin
      fu_valid <= _GEN_25;
    end
    if (reset) begin
      fu_in_wb_v <= 1'h0;
    end else if (_T) begin
      fu_in_wb_v <= io_fu_in_bits_wb_v;
    end
    if (reset) begin
      fu_in_wb_id <= 8'h0;
    end else if (_T) begin
      fu_in_wb_id <= io_fu_in_bits_wb_id;
    end
    if (reset) begin
      fu_in_wb_pc <= 32'h0;
    end else if (_T) begin
      fu_in_wb_pc <= io_fu_in_bits_wb_pc;
    end
    if (reset) begin
      fu_in_wb_instr_op <= 6'h0;
    end else if (_T) begin
      fu_in_wb_instr_op <= io_fu_in_bits_wb_instr_op;
    end
    if (reset) begin
      fu_in_wb_instr_rs_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rs_idx <= io_fu_in_bits_wb_instr_rs_idx;
    end
    if (reset) begin
      fu_in_wb_instr_rt_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rt_idx <= io_fu_in_bits_wb_instr_rt_idx;
    end
    if (reset) begin
      fu_in_wb_instr_rd_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rd_idx <= io_fu_in_bits_wb_instr_rd_idx;
    end
    if (reset) begin
      fu_in_wb_instr_shamt <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_shamt <= io_fu_in_bits_wb_instr_shamt;
    end
    if (reset) begin
      fu_in_wb_instr_func <= 6'h0;
    end else if (_T) begin
      fu_in_wb_instr_func <= io_fu_in_bits_wb_instr_func;
    end
    if (reset) begin
      fu_in_wb_rd_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_rd_idx <= io_fu_in_bits_wb_rd_idx;
    end
    if (reset) begin
      fu_in_wb_wen <= 1'h0;
    end else if (_T) begin
      fu_in_wb_wen <= io_fu_in_bits_wb_wen;
    end
    if (reset) begin
      fu_in_wb_data <= 32'h0;
    end else if (_T) begin
      fu_in_wb_data <= io_fu_in_bits_wb_data;
    end
    if (reset) begin
      fu_in_wb_is_ds <= 1'h0;
    end else if (_T) begin
      fu_in_wb_is_ds <= io_fu_in_bits_wb_is_ds;
    end
    if (reset) begin
      fu_in_wb_is_br <= 1'h0;
    end else if (_T) begin
      fu_in_wb_is_br <= io_fu_in_bits_wb_is_br;
    end
    if (reset) begin
      fu_in_wb_npc <= 32'h0;
    end else if (_T) begin
      fu_in_wb_npc <= io_fu_in_bits_wb_npc;
    end
    if (reset) begin
      fu_in_ops_fu_type <= 3'h0;
    end else if (_T) begin
      fu_in_ops_fu_type <= io_fu_in_bits_ops_fu_type;
    end
    if (reset) begin
      fu_in_ops_fu_op <= 5'h0;
    end else if (_T) begin
      fu_in_ops_fu_op <= io_fu_in_bits_ops_fu_op;
    end
    if (reset) begin
      fu_in_ops_op1 <= 32'h0;
    end else if (_T) begin
      fu_in_ops_op1 <= io_fu_in_bits_ops_op1;
    end
    if (reset) begin
      fu_in_ops_op2 <= 32'h0;
    end else if (_T) begin
      fu_in_ops_op2 <= io_fu_in_bits_ops_op2;
    end
    if (reset) begin
      fu_in_is_cached <= 1'h0;
    end else begin
      fu_in_is_cached <= _GEN_4;
    end
    if (reset) begin
      fu_in_ex_et <= 5'h0;
    end else if (_T) begin
      fu_in_ex_et <= io_fu_in_bits_ex_et;
    end
    if (reset) begin
      fu_in_ex_code <= 5'h0;
    end else if (_T) begin
      fu_in_ex_code <= io_fu_in_bits_ex_code;
    end
    if (reset) begin
      fu_in_ex_addr <= 32'h0;
    end else if (_T) begin
      fu_in_ex_addr <= io_fu_in_bits_ex_addr;
    end
    if (reset) begin
      fu_in_ex_asid <= 8'h0;
    end else if (_T) begin
      fu_in_ex_asid <= io_fu_in_bits_ex_asid;
    end
  end
endmodule
module CP0(
  input         clock,
  input         reset,
  input  [31:0] io_rport_addr,
  output [31:0] io_rport_data,
  input         io_wport_valid,
  input  [31:0] io_wport_bits_addr,
  input  [31:0] io_wport_bits_data,
  output [4:0]  io_tlbr_port_index_index,
  output [15:0] io_tlbr_port_pagemask_mask,
  output [18:0] io_tlbr_port_entry_hi_vpn,
  output [7:0]  io_tlbr_port_entry_hi_asid,
  output [19:0] io_tlbr_port_entry_lo0_pfn,
  output [2:0]  io_tlbr_port_entry_lo0_c,
  output        io_tlbr_port_entry_lo0_d,
  output        io_tlbr_port_entry_lo0_v,
  output        io_tlbr_port_entry_lo0_g,
  output [19:0] io_tlbr_port_entry_lo1_pfn,
  output [2:0]  io_tlbr_port_entry_lo1_c,
  output        io_tlbr_port_entry_lo1_d,
  output        io_tlbr_port_entry_lo1_v,
  output        io_tlbr_port_entry_lo1_g,
  input         io_tlbw_port_valid,
  input  [15:0] io_tlbw_port_bits_pagemask_mask,
  input  [18:0] io_tlbw_port_bits_entry_hi_vpn,
  input  [7:0]  io_tlbw_port_bits_entry_hi_asid,
  input  [19:0] io_tlbw_port_bits_entry_lo0_pfn,
  input  [2:0]  io_tlbw_port_bits_entry_lo0_c,
  input         io_tlbw_port_bits_entry_lo0_d,
  input         io_tlbw_port_bits_entry_lo0_v,
  input         io_tlbw_port_bits_entry_lo0_g,
  input  [19:0] io_tlbw_port_bits_entry_lo1_pfn,
  input  [2:0]  io_tlbw_port_bits_entry_lo1_c,
  input         io_tlbw_port_bits_entry_lo1_d,
  input         io_tlbw_port_bits_entry_lo1_v,
  input         io_tlbw_port_bits_entry_lo1_g,
  input         io_tlbp_port_valid,
  input         io_tlbp_port_bits_index_p,
  input  [4:0]  io_tlbp_port_bits_index_index,
  output        io_status_ERL,
  input         io_ehu_valid,
  output        io_ehu_ip7,
  input  [4:0]  io_ehu_ex_et,
  input  [4:0]  io_ehu_ex_code,
  input  [31:0] io_ehu_ex_addr,
  input  [7:0]  io_ehu_ex_asid,
  input  [31:0] io_ehu_wb_pc,
  input         io_ehu_wb_is_ds,
  input         io_ehu_wb_is_br,
  input  [31:0] io_ehu_wb_npc,
  output        io_ex_flush_valid,
  output [31:0] io_ex_flush_bits_br_target
);
  reg  cpr_index_p; // @[cp0.scala 12:26]
  reg [31:0] _RAND_0;
  reg [4:0] cpr_index_index; // @[cp0.scala 12:26]
  reg [31:0] _RAND_1;
  reg [19:0] cpr_entry_lo0_pfn; // @[cp0.scala 13:26]
  reg [31:0] _RAND_2;
  reg [2:0] cpr_entry_lo0_c; // @[cp0.scala 13:26]
  reg [31:0] _RAND_3;
  reg  cpr_entry_lo0_d; // @[cp0.scala 13:26]
  reg [31:0] _RAND_4;
  reg  cpr_entry_lo0_v; // @[cp0.scala 13:26]
  reg [31:0] _RAND_5;
  reg  cpr_entry_lo0_g; // @[cp0.scala 13:26]
  reg [31:0] _RAND_6;
  reg [19:0] cpr_entry_lo1_pfn; // @[cp0.scala 14:26]
  reg [31:0] _RAND_7;
  reg [2:0] cpr_entry_lo1_c; // @[cp0.scala 14:26]
  reg [31:0] _RAND_8;
  reg  cpr_entry_lo1_d; // @[cp0.scala 14:26]
  reg [31:0] _RAND_9;
  reg  cpr_entry_lo1_v; // @[cp0.scala 14:26]
  reg [31:0] _RAND_10;
  reg  cpr_entry_lo1_g; // @[cp0.scala 14:26]
  reg [31:0] _RAND_11;
  reg [8:0] cpr_context_ptebase; // @[cp0.scala 15:26]
  reg [31:0] _RAND_12;
  reg [18:0] cpr_context_badvpn2; // @[cp0.scala 15:26]
  reg [31:0] _RAND_13;
  reg [15:0] cpr_pagemask_mask; // @[cp0.scala 16:26]
  reg [31:0] _RAND_14;
  reg [4:0] cpr_wired_bound; // @[cp0.scala 17:26]
  reg [31:0] _RAND_15;
  reg [31:0] cpr_badvaddr; // @[cp0.scala 19:30]
  reg [31:0] _RAND_16;
  reg [31:0] cpr_count; // @[cp0.scala 20:30]
  reg [31:0] _RAND_17;
  reg [18:0] cpr_entry_hi_vpn; // @[cp0.scala 21:26]
  reg [31:0] _RAND_18;
  reg [7:0] cpr_entry_hi_asid; // @[cp0.scala 21:26]
  reg [31:0] _RAND_19;
  reg [31:0] cpr_compare; // @[cp0.scala 22:30]
  reg [31:0] _RAND_20;
  reg [3:0] cpr_status_CU; // @[cp0.scala 23:26]
  reg [31:0] _RAND_21;
  reg  cpr_status_RP; // @[cp0.scala 23:26]
  reg [31:0] _RAND_22;
  reg  cpr_status_RE; // @[cp0.scala 23:26]
  reg [31:0] _RAND_23;
  reg  cpr_status_BEV; // @[cp0.scala 23:26]
  reg [31:0] _RAND_24;
  reg  cpr_status_TS; // @[cp0.scala 23:26]
  reg [31:0] _RAND_25;
  reg  cpr_status_SR; // @[cp0.scala 23:26]
  reg [31:0] _RAND_26;
  reg  cpr_status_NMI; // @[cp0.scala 23:26]
  reg [31:0] _RAND_27;
  reg  cpr_status_IM_0; // @[cp0.scala 23:26]
  reg [31:0] _RAND_28;
  reg  cpr_status_IM_1; // @[cp0.scala 23:26]
  reg [31:0] _RAND_29;
  reg  cpr_status_IM_2; // @[cp0.scala 23:26]
  reg [31:0] _RAND_30;
  reg  cpr_status_IM_3; // @[cp0.scala 23:26]
  reg [31:0] _RAND_31;
  reg  cpr_status_IM_4; // @[cp0.scala 23:26]
  reg [31:0] _RAND_32;
  reg  cpr_status_IM_5; // @[cp0.scala 23:26]
  reg [31:0] _RAND_33;
  reg  cpr_status_IM_6; // @[cp0.scala 23:26]
  reg [31:0] _RAND_34;
  reg  cpr_status_IM_7; // @[cp0.scala 23:26]
  reg [31:0] _RAND_35;
  reg  cpr_status_UM; // @[cp0.scala 23:26]
  reg [31:0] _RAND_36;
  reg  cpr_status_ERL; // @[cp0.scala 23:26]
  reg [31:0] _RAND_37;
  reg  cpr_status_EXL; // @[cp0.scala 23:26]
  reg [31:0] _RAND_38;
  reg  cpr_status_IE; // @[cp0.scala 23:26]
  reg [31:0] _RAND_39;
  reg  cpr_cause_BD; // @[cp0.scala 24:26]
  reg [31:0] _RAND_40;
  reg  cpr_cause_IV; // @[cp0.scala 24:26]
  reg [31:0] _RAND_41;
  reg  cpr_cause_WP; // @[cp0.scala 24:26]
  reg [31:0] _RAND_42;
  reg  cpr_cause_IP_0; // @[cp0.scala 24:26]
  reg [31:0] _RAND_43;
  reg  cpr_cause_IP_1; // @[cp0.scala 24:26]
  reg [31:0] _RAND_44;
  reg  cpr_cause_IP_7; // @[cp0.scala 24:26]
  reg [31:0] _RAND_45;
  reg [4:0] cpr_cause_ExcCode; // @[cp0.scala 24:26]
  reg [31:0] _RAND_46;
  reg [31:0] cpr_epc; // @[cp0.scala 25:30]
  reg [31:0] _RAND_47;
  reg [31:0] cpr_ebase; // @[cp0.scala 27:30]
  reg [31:0] _RAND_48;
  wire [7:0] _GEN_3 = reset ? 8'h0 : cpr_entry_hi_asid; // @[cp0.scala 30:22]
  wire [18:0] _GEN_5 = reset ? 19'h0 : cpr_entry_hi_vpn; // @[cp0.scala 30:22]
  wire [8:0] _GEN_22 = reset ? 9'h0 : cpr_context_ptebase; // @[cp0.scala 30:22]
  wire [15:0] _GEN_24 = reset ? 16'h0 : cpr_pagemask_mask; // @[cp0.scala 30:22]
  wire [4:0] _GEN_26 = reset ? 5'h0 : cpr_wired_bound; // @[cp0.scala 30:22]
  wire [3:0] _GEN_28 = reset ? 4'h1 : cpr_status_CU; // @[cp0.scala 30:22]
  wire  _GEN_29 = reset ? 1'h0 : cpr_status_RP; // @[cp0.scala 30:22]
  wire  _GEN_31 = reset ? 1'h0 : cpr_status_RE; // @[cp0.scala 30:22]
  wire  _GEN_34 = reset | cpr_status_BEV; // @[cp0.scala 30:22]
  wire  _GEN_35 = reset ? 1'h0 : cpr_status_TS; // @[cp0.scala 30:22]
  wire  _GEN_36 = reset ? 1'h0 : cpr_status_SR; // @[cp0.scala 30:22]
  wire  _GEN_37 = reset ? 1'h0 : cpr_status_NMI; // @[cp0.scala 30:22]
  wire  _GEN_40 = reset ? 1'h0 : cpr_status_IM_0; // @[cp0.scala 30:22]
  wire  _GEN_41 = reset ? 1'h0 : cpr_status_IM_1; // @[cp0.scala 30:22]
  wire  _GEN_42 = reset ? 1'h0 : cpr_status_IM_2; // @[cp0.scala 30:22]
  wire  _GEN_43 = reset ? 1'h0 : cpr_status_IM_3; // @[cp0.scala 30:22]
  wire  _GEN_44 = reset ? 1'h0 : cpr_status_IM_4; // @[cp0.scala 30:22]
  wire  _GEN_45 = reset ? 1'h0 : cpr_status_IM_5; // @[cp0.scala 30:22]
  wire  _GEN_46 = reset ? 1'h0 : cpr_status_IM_6; // @[cp0.scala 30:22]
  wire  _GEN_47 = reset ? 1'h0 : cpr_status_IM_7; // @[cp0.scala 30:22]
  wire  _GEN_51 = reset ? 1'h0 : cpr_status_UM; // @[cp0.scala 30:22]
  wire  _GEN_53 = reset ? 1'h0 : cpr_status_ERL; // @[cp0.scala 30:22]
  wire  _GEN_54 = reset ? 1'h0 : cpr_status_EXL; // @[cp0.scala 30:22]
  wire  _GEN_55 = reset ? 1'h0 : cpr_status_IE; // @[cp0.scala 30:22]
  wire  _GEN_59 = reset ? 1'h0 : cpr_cause_IP_0; // @[cp0.scala 30:22]
  wire  _GEN_60 = reset ? 1'h0 : cpr_cause_IP_1; // @[cp0.scala 30:22]
  wire  _GEN_66 = reset ? 1'h0 : cpr_cause_IP_7; // @[cp0.scala 30:22]
  wire  _GEN_68 = reset ? 1'h0 : cpr_cause_WP; // @[cp0.scala 30:22]
  wire  _GEN_69 = reset ? 1'h0 : cpr_cause_IV; // @[cp0.scala 30:22]
  wire [31:0] _T_12 = cpr_count + 32'h1; // @[cp0.scala 44:26]
  wire [31:0] _T_44 = {cpr_index_p,26'h0,cpr_index_index}; // @[cp0.scala 65:32]
  wire [31:0] _T_50 = {6'h0,cpr_entry_lo0_pfn,cpr_entry_lo0_c,cpr_entry_lo0_d,cpr_entry_lo0_v,cpr_entry_lo0_g}; // @[cp0.scala 66:36]
  wire [31:0] _T_56 = {6'h0,cpr_entry_lo1_pfn,cpr_entry_lo1_c,cpr_entry_lo1_d,cpr_entry_lo1_v,cpr_entry_lo1_g}; // @[cp0.scala 67:36]
  wire [31:0] _T_58 = {cpr_context_ptebase,cpr_context_badvpn2,4'h0}; // @[cp0.scala 68:34]
  wire [31:0] _T_60 = {3'h0,cpr_pagemask_mask,13'h0}; // @[cp0.scala 69:35]
  wire [31:0] _T_61 = {27'h0,cpr_wired_bound}; // @[cp0.scala 70:32]
  wire [31:0] _T_63 = {cpr_entry_hi_vpn,5'h0,cpr_entry_hi_asid}; // @[cp0.scala 73:35]
  wire [6:0] _T_69 = {2'h0,cpr_status_UM,1'h0,cpr_status_ERL,cpr_status_EXL,cpr_status_IE}; // @[cp0.scala 75:33]
  wire [13:0] _T_76 = {cpr_status_IM_5,cpr_status_IM_4,cpr_status_IM_3,cpr_status_IM_2,cpr_status_IM_1,cpr_status_IM_0,1'h0,_T_69}; // @[cp0.scala 75:33]
  wire [7:0] _T_82 = {cpr_status_TS,cpr_status_SR,cpr_status_NMI,1'h0,2'h0,cpr_status_IM_7,cpr_status_IM_6}; // @[cp0.scala 75:33]
  wire [31:0] _T_90 = {cpr_status_CU,cpr_status_RP,1'h0,cpr_status_RE,2'h0,cpr_status_BEV,_T_82,_T_76}; // @[cp0.scala 75:33]
  wire [13:0] _T_98 = {3'h0,1'h0,cpr_cause_IP_1,cpr_cause_IP_0,1'h0,cpr_cause_ExcCode,2'h0}; // @[cp0.scala 76:32]
  wire [31:0] _T_107 = {cpr_cause_BD,1'h0,2'h0,4'h0,cpr_cause_IV,cpr_cause_WP,6'h0,cpr_cause_IP_7,1'h0,_T_98}; // @[cp0.scala 76:32]
  wire  _T_132 = 32'h81 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_133 = _T_132 ? 32'h3e9b4d80 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_134 = 32'h80 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_135 = _T_134 ? 32'h80000080 : _T_133; // @[Mux.scala 68:16]
  wire  _T_136 = 32'h79 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_137 = _T_136 ? cpr_ebase : _T_135; // @[Mux.scala 68:16]
  wire  _T_138 = 32'h78 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_139 = _T_138 ? 32'h18000 : _T_137; // @[Mux.scala 68:16]
  wire  _T_140 = 32'h70 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_141 = _T_140 ? cpr_epc : _T_139; // @[Mux.scala 68:16]
  wire  _T_142 = 32'h68 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_143 = _T_142 ? _T_107 : _T_141; // @[Mux.scala 68:16]
  wire  _T_144 = 32'h60 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_145 = _T_144 ? _T_90 : _T_143; // @[Mux.scala 68:16]
  wire  _T_146 = 32'h58 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_147 = _T_146 ? cpr_compare : _T_145; // @[Mux.scala 68:16]
  wire  _T_148 = 32'h50 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_149 = _T_148 ? _T_63 : _T_147; // @[Mux.scala 68:16]
  wire  _T_150 = 32'h48 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_151 = _T_150 ? cpr_count : _T_149; // @[Mux.scala 68:16]
  wire  _T_152 = 32'h40 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_153 = _T_152 ? cpr_badvaddr : _T_151; // @[Mux.scala 68:16]
  wire  _T_154 = 32'h30 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_155 = _T_154 ? _T_61 : _T_153; // @[Mux.scala 68:16]
  wire  _T_156 = 32'h28 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_157 = _T_156 ? _T_60 : _T_155; // @[Mux.scala 68:16]
  wire  _T_158 = 32'h20 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_159 = _T_158 ? _T_58 : _T_157; // @[Mux.scala 68:16]
  wire  _T_160 = 32'h18 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_161 = _T_160 ? _T_56 : _T_159; // @[Mux.scala 68:16]
  wire  _T_162 = 32'h10 == io_rport_addr; // @[Mux.scala 68:19]
  wire [31:0] _T_163 = _T_162 ? _T_50 : _T_161; // @[Mux.scala 68:16]
  wire  _T_164 = 32'h0 == io_rport_addr; // @[Mux.scala 68:19]
  wire  _T_166 = ~io_ex_flush_valid; // @[cp0.scala 85:27]
  wire  _T_167 = io_wport_valid & _T_166; // @[cp0.scala 85:24]
  wire  _T_168 = 32'h0 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_174 = 32'h10 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_184 = 32'h18 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_194 = 32'h20 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_200 = 32'h28 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_206 = 32'h30 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_211 = 32'h40 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_212 = 32'h48 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_213 = 32'h50 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_219 = 32'h58 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_220 = 32'h60 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_251 = 32'h68 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_272 = 32'h70 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_273 = 32'h78 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _T_274 = 32'h79 == io_wport_bits_addr; // @[Conditional.scala 37:30]
  wire  _GEN_137 = _T_219 ? 1'h0 : _GEN_66; // @[Conditional.scala 39:67]
  wire  _GEN_166 = _T_213 ? _GEN_66 : _GEN_137; // @[Conditional.scala 39:67]
  wire  _GEN_195 = _T_212 ? _GEN_66 : _GEN_166; // @[Conditional.scala 39:67]
  wire  _GEN_225 = _T_211 ? _GEN_66 : _GEN_195; // @[Conditional.scala 39:67]
  wire  _GEN_256 = _T_206 ? _GEN_66 : _GEN_225; // @[Conditional.scala 39:67]
  wire  _GEN_288 = _T_200 ? _GEN_66 : _GEN_256; // @[Conditional.scala 39:67]
  wire  _GEN_321 = _T_194 ? _GEN_66 : _GEN_288; // @[Conditional.scala 39:67]
  wire  _GEN_359 = _T_184 ? _GEN_66 : _GEN_321; // @[Conditional.scala 39:67]
  wire  _GEN_402 = _T_174 ? _GEN_66 : _GEN_359; // @[Conditional.scala 39:67]
  wire  _GEN_446 = _T_168 ? _GEN_66 : _GEN_402; // @[Conditional.scala 40:58]
  wire  _GEN_490 = _T_167 ? _GEN_446 : _GEN_66; // @[cp0.scala 85:47]
  wire  _T_278 = io_tlbw_port_valid & _T_166; // @[cp0.scala 116:28]
  wire [31:0] _T_280 = {3'h0,io_tlbw_port_bits_pagemask_mask,13'h0}; // @[cp0.scala 118:39]
  wire [31:0] _T_287 = {io_tlbw_port_bits_entry_hi_vpn,5'h0,io_tlbw_port_bits_entry_hi_asid}; // @[cp0.scala 119:39]
  wire [31:0] _T_298 = {6'h0,io_tlbw_port_bits_entry_lo0_pfn,io_tlbw_port_bits_entry_lo0_c,io_tlbw_port_bits_entry_lo0_d,io_tlbw_port_bits_entry_lo0_v,io_tlbw_port_bits_entry_lo0_g}; // @[cp0.scala 120:41]
  wire [31:0] _T_313 = {6'h0,io_tlbw_port_bits_entry_lo1_pfn,io_tlbw_port_bits_entry_lo1_c,io_tlbw_port_bits_entry_lo1_d,io_tlbw_port_bits_entry_lo1_v,io_tlbw_port_bits_entry_lo1_g}; // @[cp0.scala 121:41]
  wire  _T_324 = io_tlbp_port_valid & _T_166; // @[cp0.scala 124:28]
  wire  _T_326 = ~io_tlbp_port_bits_index_p; // @[cp0.scala 126:11]
  wire  _T_328 = ~cpr_status_ERL; // @[cp0.scala 133:21]
  wire  _T_329 = ~cpr_status_EXL; // @[cp0.scala 133:40]
  wire  _T_330 = _T_328 & _T_329; // @[cp0.scala 133:37]
  wire  intr_enable = _T_330 & cpr_status_IE; // @[cp0.scala 133:56]
  wire [7:0] _T_337 = {cpr_cause_IP_7,1'h0,2'h0,2'h0,cpr_cause_IP_1,cpr_cause_IP_0}; // @[cp0.scala 134:34]
  wire [7:0] _T_344 = {cpr_status_IM_7,cpr_status_IM_6,cpr_status_IM_5,cpr_status_IM_4,cpr_status_IM_3,cpr_status_IM_2,cpr_status_IM_1,cpr_status_IM_0}; // @[cp0.scala 134:57]
  wire [7:0] _T_345 = _T_337 & _T_344; // @[cp0.scala 134:41]
  wire  _T_346 = _T_345 != 8'h0; // @[cp0.scala 134:65]
  wire  intr_valid = _T_346 & intr_enable; // @[cp0.scala 134:69]
  wire  intr_flush = io_ehu_valid & intr_valid; // @[cp0.scala 135:33]
  wire  _T_347 = io_ehu_ex_et != 5'h0; // @[cp0.scala 136:47]
  wire  ex_flush = io_ehu_valid & _T_347; // @[cp0.scala 136:31]
  wire  _T_348 = ~ex_flush; // @[cp0.scala 137:34]
  wire  is_intr_ex = intr_flush & _T_348; // @[cp0.scala 137:31]
  wire  _T_350 = io_ehu_ex_et != 5'h16; // @[cp0.scala 141:24]
  wire  _T_353 = is_intr_ex & io_ehu_wb_is_br; // @[cp0.scala 147:23]
  wire  _T_354 = ~io_ehu_wb_is_br; // @[cp0.scala 148:26]
  wire  _T_355 = is_intr_ex & _T_354; // @[cp0.scala 148:23]
  wire [31:0] _T_357 = io_ehu_wb_pc - 32'h4; // @[cp0.scala 149:34]
  wire  _T_361 = io_ehu_ex_et == 5'h0; // @[cp0.scala 152:45]
  wire  _T_365 = io_ehu_ex_et == 5'h16; // @[cp0.scala 158:31]
  wire  _T_366 = io_ehu_ex_et == 5'h6; // @[cp0.scala 162:24]
  wire  _T_367 = io_ehu_ex_et == 5'h8; // @[cp0.scala 164:30]
  wire  _T_368 = io_ehu_ex_et == 5'h9; // @[cp0.scala 165:20]
  wire  _T_369 = _T_367 | _T_368; // @[cp0.scala 164:45]
  wire  _T_370 = io_ehu_ex_et == 5'h7; // @[cp0.scala 166:20]
  wire  _T_371 = _T_369 | _T_370; // @[cp0.scala 165:35]
  wire  _T_374 = io_ehu_ex_et != 5'h7; // @[cp0.scala 170:26]
  wire  _T_377 = is_intr_ex & cpr_cause_IV; // @[cp0.scala 178:17]
  wire [9:0] _T_378 = _T_377 ? 10'h200 : 10'h180; // @[Mux.scala 87:16]
  wire [9:0] _T_379 = _T_370 ? 10'h0 : _T_378; // @[Mux.scala 87:16]
  wire [9:0] offset = cpr_status_EXL ? 10'h180 : _T_379; // @[Mux.scala 87:16]
  wire [31:0] _GEN_559 = {{22'd0}, offset}; // @[cp0.scala 181:47]
  wire [31:0] _T_383 = 32'hbfc00200 + _GEN_559; // @[cp0.scala 181:47]
  wire [31:0] _T_385 = 32'h80000000 + _GEN_559; // @[cp0.scala 182:21]
  wire [31:0] _T_386 = cpr_status_BEV ? _T_383 : _T_385; // @[cp0.scala 181:8]
  wire  _T_388 = cpr_compare == cpr_count; // @[cp0.scala 184:21]
  assign io_rport_data = _T_164 ? _T_44 : _T_163; // @[cp0.scala 64:17]
  assign io_tlbr_port_index_index = cpr_index_index; // @[cp0.scala 111:22]
  assign io_tlbr_port_pagemask_mask = cpr_pagemask_mask; // @[cp0.scala 110:25]
  assign io_tlbr_port_entry_hi_vpn = cpr_entry_hi_vpn; // @[cp0.scala 112:25]
  assign io_tlbr_port_entry_hi_asid = cpr_entry_hi_asid; // @[cp0.scala 112:25]
  assign io_tlbr_port_entry_lo0_pfn = cpr_entry_lo0_pfn; // @[cp0.scala 113:26]
  assign io_tlbr_port_entry_lo0_c = cpr_entry_lo0_c; // @[cp0.scala 113:26]
  assign io_tlbr_port_entry_lo0_d = cpr_entry_lo0_d; // @[cp0.scala 113:26]
  assign io_tlbr_port_entry_lo0_v = cpr_entry_lo0_v; // @[cp0.scala 113:26]
  assign io_tlbr_port_entry_lo0_g = cpr_entry_lo0_g; // @[cp0.scala 113:26]
  assign io_tlbr_port_entry_lo1_pfn = cpr_entry_lo1_pfn; // @[cp0.scala 114:26]
  assign io_tlbr_port_entry_lo1_c = cpr_entry_lo1_c; // @[cp0.scala 114:26]
  assign io_tlbr_port_entry_lo1_d = cpr_entry_lo1_d; // @[cp0.scala 114:26]
  assign io_tlbr_port_entry_lo1_v = cpr_entry_lo1_v; // @[cp0.scala 114:26]
  assign io_tlbr_port_entry_lo1_g = cpr_entry_lo1_g; // @[cp0.scala 114:26]
  assign io_status_ERL = cpr_status_ERL; // @[cp0.scala 60:13]
  assign io_ehu_ip7 = cpr_cause_IP_7; // @[cp0.scala 138:14]
  assign io_ex_flush_valid = intr_flush | ex_flush; // @[cp0.scala 139:21]
  assign io_ex_flush_bits_br_target = _T_365 ? cpr_epc : _T_386; // @[cp0.scala 179:30]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cpr_index_p = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cpr_index_index = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cpr_entry_lo0_pfn = _RAND_2[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cpr_entry_lo0_c = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  cpr_entry_lo0_d = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  cpr_entry_lo0_v = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  cpr_entry_lo0_g = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  cpr_entry_lo1_pfn = _RAND_7[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  cpr_entry_lo1_c = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  cpr_entry_lo1_d = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  cpr_entry_lo1_v = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  cpr_entry_lo1_g = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  cpr_context_ptebase = _RAND_12[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  cpr_context_badvpn2 = _RAND_13[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  cpr_pagemask_mask = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  cpr_wired_bound = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  cpr_badvaddr = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  cpr_count = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  cpr_entry_hi_vpn = _RAND_18[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  cpr_entry_hi_asid = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  cpr_compare = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  cpr_status_CU = _RAND_21[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  cpr_status_RP = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  cpr_status_RE = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  cpr_status_BEV = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  cpr_status_TS = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  cpr_status_SR = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  cpr_status_NMI = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  cpr_status_IM_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  cpr_status_IM_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  cpr_status_IM_2 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  cpr_status_IM_3 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  cpr_status_IM_4 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  cpr_status_IM_5 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  cpr_status_IM_6 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  cpr_status_IM_7 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  cpr_status_UM = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  cpr_status_ERL = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  cpr_status_EXL = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  cpr_status_IE = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  cpr_cause_BD = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  cpr_cause_IV = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  cpr_cause_WP = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  cpr_cause_IP_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  cpr_cause_IP_1 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  cpr_cause_IP_7 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  cpr_cause_ExcCode = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  cpr_epc = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  cpr_ebase = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T_324) begin
      cpr_index_p <= io_tlbp_port_bits_index_p;
    end else if (reset) begin
      cpr_index_p <= 1'h0;
    end
    if (_T_324) begin
      if (_T_326) begin
        cpr_index_index <= io_tlbp_port_bits_index_index;
      end else if (_T_167) begin
        if (_T_168) begin
          cpr_index_index <= io_wport_bits_data[4:0];
        end else if (reset) begin
          cpr_index_index <= 5'h0;
        end
      end else if (reset) begin
        cpr_index_index <= 5'h0;
      end
    end else if (_T_167) begin
      if (_T_168) begin
        cpr_index_index <= io_wport_bits_data[4:0];
      end else if (reset) begin
        cpr_index_index <= 5'h0;
      end
    end else if (reset) begin
      cpr_index_index <= 5'h0;
    end
    if (_T_278) begin
      cpr_entry_lo0_pfn <= _T_298[25:6];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo0_pfn <= 20'h0;
        end
      end else if (_T_174) begin
        cpr_entry_lo0_pfn <= io_wport_bits_data[25:6];
      end else if (reset) begin
        cpr_entry_lo0_pfn <= 20'h0;
      end
    end else if (reset) begin
      cpr_entry_lo0_pfn <= 20'h0;
    end
    if (_T_278) begin
      cpr_entry_lo0_c <= _T_298[5:3];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo0_c <= 3'h0;
        end
      end else if (_T_174) begin
        cpr_entry_lo0_c <= io_wport_bits_data[5:3];
      end else if (reset) begin
        cpr_entry_lo0_c <= 3'h0;
      end
    end else if (reset) begin
      cpr_entry_lo0_c <= 3'h0;
    end
    if (_T_278) begin
      cpr_entry_lo0_d <= _T_298[2];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo0_d <= 1'h0;
        end
      end else if (_T_174) begin
        cpr_entry_lo0_d <= io_wport_bits_data[2];
      end else if (reset) begin
        cpr_entry_lo0_d <= 1'h0;
      end
    end else if (reset) begin
      cpr_entry_lo0_d <= 1'h0;
    end
    if (_T_278) begin
      cpr_entry_lo0_v <= _T_298[1];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo0_v <= 1'h0;
        end
      end else if (_T_174) begin
        cpr_entry_lo0_v <= io_wport_bits_data[1];
      end else if (reset) begin
        cpr_entry_lo0_v <= 1'h0;
      end
    end else if (reset) begin
      cpr_entry_lo0_v <= 1'h0;
    end
    if (_T_278) begin
      cpr_entry_lo0_g <= _T_298[0];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo0_g <= 1'h0;
        end
      end else if (_T_174) begin
        cpr_entry_lo0_g <= io_wport_bits_data[0];
      end else if (reset) begin
        cpr_entry_lo0_g <= 1'h0;
      end
    end else if (reset) begin
      cpr_entry_lo0_g <= 1'h0;
    end
    if (_T_278) begin
      cpr_entry_lo1_pfn <= _T_313[25:6];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo1_pfn <= 20'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_entry_lo1_pfn <= 20'h0;
        end
      end else if (_T_184) begin
        cpr_entry_lo1_pfn <= io_wport_bits_data[25:6];
      end else if (reset) begin
        cpr_entry_lo1_pfn <= 20'h0;
      end
    end else if (reset) begin
      cpr_entry_lo1_pfn <= 20'h0;
    end
    if (_T_278) begin
      cpr_entry_lo1_c <= _T_313[5:3];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo1_c <= 3'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_entry_lo1_c <= 3'h0;
        end
      end else if (_T_184) begin
        cpr_entry_lo1_c <= io_wport_bits_data[5:3];
      end else if (reset) begin
        cpr_entry_lo1_c <= 3'h0;
      end
    end else if (reset) begin
      cpr_entry_lo1_c <= 3'h0;
    end
    if (_T_278) begin
      cpr_entry_lo1_d <= _T_313[2];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo1_d <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_entry_lo1_d <= 1'h0;
        end
      end else if (_T_184) begin
        cpr_entry_lo1_d <= io_wport_bits_data[2];
      end else if (reset) begin
        cpr_entry_lo1_d <= 1'h0;
      end
    end else if (reset) begin
      cpr_entry_lo1_d <= 1'h0;
    end
    if (_T_278) begin
      cpr_entry_lo1_v <= _T_313[1];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo1_v <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_entry_lo1_v <= 1'h0;
        end
      end else if (_T_184) begin
        cpr_entry_lo1_v <= io_wport_bits_data[1];
      end else if (reset) begin
        cpr_entry_lo1_v <= 1'h0;
      end
    end else if (reset) begin
      cpr_entry_lo1_v <= 1'h0;
    end
    if (_T_278) begin
      cpr_entry_lo1_g <= _T_313[0];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_entry_lo1_g <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_entry_lo1_g <= 1'h0;
        end
      end else if (_T_184) begin
        cpr_entry_lo1_g <= io_wport_bits_data[0];
      end else if (reset) begin
        cpr_entry_lo1_g <= 1'h0;
      end
    end else if (reset) begin
      cpr_entry_lo1_g <= 1'h0;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_context_ptebase <= 9'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_context_ptebase <= 9'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_context_ptebase <= 9'h0;
        end
      end else if (_T_194) begin
        cpr_context_ptebase <= io_wport_bits_data[31:23];
      end else if (reset) begin
        cpr_context_ptebase <= 9'h0;
      end
    end else begin
      cpr_context_ptebase <= _GEN_22;
    end
    if (io_ex_flush_valid) begin
      if (_T_366) begin
        if (reset) begin
          cpr_context_badvpn2 <= 19'h0;
        end
      end else if (_T_371) begin
        cpr_context_badvpn2 <= io_ehu_ex_addr[31:13];
      end else if (reset) begin
        cpr_context_badvpn2 <= 19'h0;
      end
    end else if (reset) begin
      cpr_context_badvpn2 <= 19'h0;
    end
    if (_T_278) begin
      cpr_pagemask_mask <= _T_280[28:13];
    end else if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_pagemask_mask <= 16'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_pagemask_mask <= 16'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_pagemask_mask <= 16'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_pagemask_mask <= 16'h0;
        end
      end else if (_T_200) begin
        cpr_pagemask_mask <= io_wport_bits_data[28:13];
      end else begin
        cpr_pagemask_mask <= _GEN_24;
      end
    end else begin
      cpr_pagemask_mask <= _GEN_24;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_wired_bound <= 5'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_wired_bound <= 5'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_wired_bound <= 5'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_wired_bound <= 5'h0;
        end
      end else if (_T_200) begin
        cpr_wired_bound <= _GEN_26;
      end else if (_T_206) begin
        cpr_wired_bound <= io_wport_bits_data[4:0];
      end else begin
        cpr_wired_bound <= _GEN_26;
      end
    end else begin
      cpr_wired_bound <= _GEN_26;
    end
    if (reset) begin
      cpr_badvaddr <= 32'h0;
    end else if (io_ex_flush_valid) begin
      if (_T_366) begin
        cpr_badvaddr <= io_ehu_ex_addr;
      end else if (_T_371) begin
        cpr_badvaddr <= io_ehu_ex_addr;
      end else if (_T_167) begin
        if (!(_T_168)) begin
          if (!(_T_174)) begin
            if (!(_T_184)) begin
              if (!(_T_194)) begin
                if (!(_T_200)) begin
                  if (!(_T_206)) begin
                    if (_T_211) begin
                      cpr_badvaddr <= io_wport_bits_data;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else if (_T_167) begin
      if (!(_T_168)) begin
        if (!(_T_174)) begin
          if (!(_T_184)) begin
            if (!(_T_194)) begin
              if (!(_T_200)) begin
                if (!(_T_206)) begin
                  if (_T_211) begin
                    cpr_badvaddr <= io_wport_bits_data;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cpr_count <= 32'h1;
    end else begin
      cpr_count <= _T_12;
    end
    if (io_ex_flush_valid) begin
      if (_T_366) begin
        if (_T_278) begin
          cpr_entry_hi_vpn <= _T_287[31:13];
        end else if (_T_167) begin
          if (_T_168) begin
            if (reset) begin
              cpr_entry_hi_vpn <= 19'h0;
            end
          end else if (_T_174) begin
            if (reset) begin
              cpr_entry_hi_vpn <= 19'h0;
            end
          end else if (_T_184) begin
            if (reset) begin
              cpr_entry_hi_vpn <= 19'h0;
            end
          end else if (_T_194) begin
            if (reset) begin
              cpr_entry_hi_vpn <= 19'h0;
            end
          end else if (_T_200) begin
            cpr_entry_hi_vpn <= _GEN_5;
          end else if (_T_206) begin
            cpr_entry_hi_vpn <= _GEN_5;
          end else if (_T_211) begin
            cpr_entry_hi_vpn <= _GEN_5;
          end else if (_T_212) begin
            cpr_entry_hi_vpn <= _GEN_5;
          end else if (_T_213) begin
            cpr_entry_hi_vpn <= io_wport_bits_data[31:13];
          end else begin
            cpr_entry_hi_vpn <= _GEN_5;
          end
        end else begin
          cpr_entry_hi_vpn <= _GEN_5;
        end
      end else if (_T_371) begin
        cpr_entry_hi_vpn <= io_ehu_ex_addr[31:13];
      end else if (_T_278) begin
        cpr_entry_hi_vpn <= _T_287[31:13];
      end else if (_T_167) begin
        if (_T_168) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_174) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_184) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_194) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_200) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_206) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_211) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_212) begin
          cpr_entry_hi_vpn <= _GEN_5;
        end else if (_T_213) begin
          cpr_entry_hi_vpn <= io_wport_bits_data[31:13];
        end else begin
          cpr_entry_hi_vpn <= _GEN_5;
        end
      end else begin
        cpr_entry_hi_vpn <= _GEN_5;
      end
    end else if (_T_278) begin
      cpr_entry_hi_vpn <= _T_287[31:13];
    end else if (_T_167) begin
      if (_T_168) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_174) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_184) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_194) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_200) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_206) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_211) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_212) begin
        cpr_entry_hi_vpn <= _GEN_5;
      end else if (_T_213) begin
        cpr_entry_hi_vpn <= io_wport_bits_data[31:13];
      end else begin
        cpr_entry_hi_vpn <= _GEN_5;
      end
    end else begin
      cpr_entry_hi_vpn <= _GEN_5;
    end
    if (io_ex_flush_valid) begin
      if (_T_366) begin
        if (_T_278) begin
          cpr_entry_hi_asid <= _T_287[7:0];
        end else if (_T_167) begin
          if (_T_168) begin
            if (reset) begin
              cpr_entry_hi_asid <= 8'h0;
            end
          end else if (_T_174) begin
            if (reset) begin
              cpr_entry_hi_asid <= 8'h0;
            end
          end else if (_T_184) begin
            if (reset) begin
              cpr_entry_hi_asid <= 8'h0;
            end
          end else if (_T_194) begin
            if (reset) begin
              cpr_entry_hi_asid <= 8'h0;
            end
          end else if (_T_200) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_206) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_211) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_212) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_213) begin
            cpr_entry_hi_asid <= io_wport_bits_data[7:0];
          end else begin
            cpr_entry_hi_asid <= _GEN_3;
          end
        end else begin
          cpr_entry_hi_asid <= _GEN_3;
        end
      end else if (_T_371) begin
        if (_T_374) begin
          cpr_entry_hi_asid <= io_ehu_ex_asid;
        end else if (_T_278) begin
          cpr_entry_hi_asid <= _T_287[7:0];
        end else if (_T_167) begin
          if (_T_168) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_174) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_184) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_194) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_200) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_206) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_211) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_212) begin
            cpr_entry_hi_asid <= _GEN_3;
          end else if (_T_213) begin
            cpr_entry_hi_asid <= io_wport_bits_data[7:0];
          end else begin
            cpr_entry_hi_asid <= _GEN_3;
          end
        end else begin
          cpr_entry_hi_asid <= _GEN_3;
        end
      end else if (_T_278) begin
        cpr_entry_hi_asid <= _T_287[7:0];
      end else if (_T_167) begin
        if (_T_168) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_174) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_184) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_194) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_200) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_206) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_211) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_212) begin
          cpr_entry_hi_asid <= _GEN_3;
        end else if (_T_213) begin
          cpr_entry_hi_asid <= io_wport_bits_data[7:0];
        end else begin
          cpr_entry_hi_asid <= _GEN_3;
        end
      end else begin
        cpr_entry_hi_asid <= _GEN_3;
      end
    end else if (_T_278) begin
      cpr_entry_hi_asid <= _T_287[7:0];
    end else if (_T_167) begin
      if (_T_168) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_174) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_184) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_194) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_200) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_206) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_211) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_212) begin
        cpr_entry_hi_asid <= _GEN_3;
      end else if (_T_213) begin
        cpr_entry_hi_asid <= io_wport_bits_data[7:0];
      end else begin
        cpr_entry_hi_asid <= _GEN_3;
      end
    end else begin
      cpr_entry_hi_asid <= _GEN_3;
    end
    if (reset) begin
      cpr_compare <= 32'hffffffff;
    end else if (_T_167) begin
      if (!(_T_168)) begin
        if (!(_T_174)) begin
          if (!(_T_184)) begin
            if (!(_T_194)) begin
              if (!(_T_200)) begin
                if (!(_T_206)) begin
                  if (!(_T_211)) begin
                    if (!(_T_212)) begin
                      if (!(_T_213)) begin
                        if (_T_219) begin
                          cpr_compare <= io_wport_bits_data;
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_CU <= 4'h1;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_CU <= 4'h1;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_CU <= 4'h1;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_CU <= 4'h1;
        end
      end else if (_T_200) begin
        cpr_status_CU <= _GEN_28;
      end else if (_T_206) begin
        cpr_status_CU <= _GEN_28;
      end else if (_T_211) begin
        cpr_status_CU <= _GEN_28;
      end else if (_T_212) begin
        cpr_status_CU <= _GEN_28;
      end else if (_T_213) begin
        cpr_status_CU <= _GEN_28;
      end else if (_T_219) begin
        cpr_status_CU <= _GEN_28;
      end else if (_T_220) begin
        cpr_status_CU <= io_wport_bits_data[31:28];
      end else begin
        cpr_status_CU <= _GEN_28;
      end
    end else begin
      cpr_status_CU <= _GEN_28;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_RP <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_RP <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_RP <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_RP <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_RP <= _GEN_29;
      end else if (_T_206) begin
        cpr_status_RP <= _GEN_29;
      end else if (_T_211) begin
        cpr_status_RP <= _GEN_29;
      end else if (_T_212) begin
        cpr_status_RP <= _GEN_29;
      end else if (_T_213) begin
        cpr_status_RP <= _GEN_29;
      end else if (_T_219) begin
        cpr_status_RP <= _GEN_29;
      end else if (_T_220) begin
        cpr_status_RP <= io_wport_bits_data[27];
      end else begin
        cpr_status_RP <= _GEN_29;
      end
    end else begin
      cpr_status_RP <= _GEN_29;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_RE <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_RE <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_RE <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_RE <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_RE <= _GEN_31;
      end else if (_T_206) begin
        cpr_status_RE <= _GEN_31;
      end else if (_T_211) begin
        cpr_status_RE <= _GEN_31;
      end else if (_T_212) begin
        cpr_status_RE <= _GEN_31;
      end else if (_T_213) begin
        cpr_status_RE <= _GEN_31;
      end else if (_T_219) begin
        cpr_status_RE <= _GEN_31;
      end else if (_T_220) begin
        cpr_status_RE <= io_wport_bits_data[25];
      end else begin
        cpr_status_RE <= _GEN_31;
      end
    end else begin
      cpr_status_RE <= _GEN_31;
    end
    if (_T_167) begin
      if (_T_168) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_174) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_184) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_194) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_200) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_206) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_211) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_212) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_213) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_219) begin
        cpr_status_BEV <= _GEN_34;
      end else if (_T_220) begin
        cpr_status_BEV <= io_wport_bits_data[22];
      end else begin
        cpr_status_BEV <= _GEN_34;
      end
    end else begin
      cpr_status_BEV <= _GEN_34;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_TS <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_TS <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_TS <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_TS <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_TS <= _GEN_35;
      end else if (_T_206) begin
        cpr_status_TS <= _GEN_35;
      end else if (_T_211) begin
        cpr_status_TS <= _GEN_35;
      end else if (_T_212) begin
        cpr_status_TS <= _GEN_35;
      end else if (_T_213) begin
        cpr_status_TS <= _GEN_35;
      end else if (_T_219) begin
        cpr_status_TS <= _GEN_35;
      end else if (_T_220) begin
        cpr_status_TS <= io_wport_bits_data[21];
      end else begin
        cpr_status_TS <= _GEN_35;
      end
    end else begin
      cpr_status_TS <= _GEN_35;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_SR <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_SR <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_SR <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_SR <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_SR <= _GEN_36;
      end else if (_T_206) begin
        cpr_status_SR <= _GEN_36;
      end else if (_T_211) begin
        cpr_status_SR <= _GEN_36;
      end else if (_T_212) begin
        cpr_status_SR <= _GEN_36;
      end else if (_T_213) begin
        cpr_status_SR <= _GEN_36;
      end else if (_T_219) begin
        cpr_status_SR <= _GEN_36;
      end else if (_T_220) begin
        cpr_status_SR <= io_wport_bits_data[20];
      end else begin
        cpr_status_SR <= _GEN_36;
      end
    end else begin
      cpr_status_SR <= _GEN_36;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_NMI <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_NMI <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_NMI <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_NMI <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_NMI <= _GEN_37;
      end else if (_T_206) begin
        cpr_status_NMI <= _GEN_37;
      end else if (_T_211) begin
        cpr_status_NMI <= _GEN_37;
      end else if (_T_212) begin
        cpr_status_NMI <= _GEN_37;
      end else if (_T_213) begin
        cpr_status_NMI <= _GEN_37;
      end else if (_T_219) begin
        cpr_status_NMI <= _GEN_37;
      end else if (_T_220) begin
        cpr_status_NMI <= io_wport_bits_data[19];
      end else begin
        cpr_status_NMI <= _GEN_37;
      end
    end else begin
      cpr_status_NMI <= _GEN_37;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_0 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_0 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_0 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_0 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_0 <= _GEN_40;
      end else if (_T_206) begin
        cpr_status_IM_0 <= _GEN_40;
      end else if (_T_211) begin
        cpr_status_IM_0 <= _GEN_40;
      end else if (_T_212) begin
        cpr_status_IM_0 <= _GEN_40;
      end else if (_T_213) begin
        cpr_status_IM_0 <= _GEN_40;
      end else if (_T_219) begin
        cpr_status_IM_0 <= _GEN_40;
      end else if (_T_220) begin
        cpr_status_IM_0 <= io_wport_bits_data[8];
      end else begin
        cpr_status_IM_0 <= _GEN_40;
      end
    end else begin
      cpr_status_IM_0 <= _GEN_40;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_1 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_1 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_1 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_1 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_1 <= _GEN_41;
      end else if (_T_206) begin
        cpr_status_IM_1 <= _GEN_41;
      end else if (_T_211) begin
        cpr_status_IM_1 <= _GEN_41;
      end else if (_T_212) begin
        cpr_status_IM_1 <= _GEN_41;
      end else if (_T_213) begin
        cpr_status_IM_1 <= _GEN_41;
      end else if (_T_219) begin
        cpr_status_IM_1 <= _GEN_41;
      end else if (_T_220) begin
        cpr_status_IM_1 <= io_wport_bits_data[9];
      end else begin
        cpr_status_IM_1 <= _GEN_41;
      end
    end else begin
      cpr_status_IM_1 <= _GEN_41;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_2 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_2 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_2 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_2 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_2 <= _GEN_42;
      end else if (_T_206) begin
        cpr_status_IM_2 <= _GEN_42;
      end else if (_T_211) begin
        cpr_status_IM_2 <= _GEN_42;
      end else if (_T_212) begin
        cpr_status_IM_2 <= _GEN_42;
      end else if (_T_213) begin
        cpr_status_IM_2 <= _GEN_42;
      end else if (_T_219) begin
        cpr_status_IM_2 <= _GEN_42;
      end else if (_T_220) begin
        cpr_status_IM_2 <= io_wport_bits_data[10];
      end else begin
        cpr_status_IM_2 <= _GEN_42;
      end
    end else begin
      cpr_status_IM_2 <= _GEN_42;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_3 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_3 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_3 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_3 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_3 <= _GEN_43;
      end else if (_T_206) begin
        cpr_status_IM_3 <= _GEN_43;
      end else if (_T_211) begin
        cpr_status_IM_3 <= _GEN_43;
      end else if (_T_212) begin
        cpr_status_IM_3 <= _GEN_43;
      end else if (_T_213) begin
        cpr_status_IM_3 <= _GEN_43;
      end else if (_T_219) begin
        cpr_status_IM_3 <= _GEN_43;
      end else if (_T_220) begin
        cpr_status_IM_3 <= io_wport_bits_data[11];
      end else begin
        cpr_status_IM_3 <= _GEN_43;
      end
    end else begin
      cpr_status_IM_3 <= _GEN_43;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_4 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_4 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_4 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_4 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_4 <= _GEN_44;
      end else if (_T_206) begin
        cpr_status_IM_4 <= _GEN_44;
      end else if (_T_211) begin
        cpr_status_IM_4 <= _GEN_44;
      end else if (_T_212) begin
        cpr_status_IM_4 <= _GEN_44;
      end else if (_T_213) begin
        cpr_status_IM_4 <= _GEN_44;
      end else if (_T_219) begin
        cpr_status_IM_4 <= _GEN_44;
      end else if (_T_220) begin
        cpr_status_IM_4 <= io_wport_bits_data[12];
      end else begin
        cpr_status_IM_4 <= _GEN_44;
      end
    end else begin
      cpr_status_IM_4 <= _GEN_44;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_5 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_5 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_5 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_5 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_5 <= _GEN_45;
      end else if (_T_206) begin
        cpr_status_IM_5 <= _GEN_45;
      end else if (_T_211) begin
        cpr_status_IM_5 <= _GEN_45;
      end else if (_T_212) begin
        cpr_status_IM_5 <= _GEN_45;
      end else if (_T_213) begin
        cpr_status_IM_5 <= _GEN_45;
      end else if (_T_219) begin
        cpr_status_IM_5 <= _GEN_45;
      end else if (_T_220) begin
        cpr_status_IM_5 <= io_wport_bits_data[13];
      end else begin
        cpr_status_IM_5 <= _GEN_45;
      end
    end else begin
      cpr_status_IM_5 <= _GEN_45;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_6 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_6 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_6 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_6 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_6 <= _GEN_46;
      end else if (_T_206) begin
        cpr_status_IM_6 <= _GEN_46;
      end else if (_T_211) begin
        cpr_status_IM_6 <= _GEN_46;
      end else if (_T_212) begin
        cpr_status_IM_6 <= _GEN_46;
      end else if (_T_213) begin
        cpr_status_IM_6 <= _GEN_46;
      end else if (_T_219) begin
        cpr_status_IM_6 <= _GEN_46;
      end else if (_T_220) begin
        cpr_status_IM_6 <= io_wport_bits_data[14];
      end else begin
        cpr_status_IM_6 <= _GEN_46;
      end
    end else begin
      cpr_status_IM_6 <= _GEN_46;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IM_7 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IM_7 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IM_7 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IM_7 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IM_7 <= _GEN_47;
      end else if (_T_206) begin
        cpr_status_IM_7 <= _GEN_47;
      end else if (_T_211) begin
        cpr_status_IM_7 <= _GEN_47;
      end else if (_T_212) begin
        cpr_status_IM_7 <= _GEN_47;
      end else if (_T_213) begin
        cpr_status_IM_7 <= _GEN_47;
      end else if (_T_219) begin
        cpr_status_IM_7 <= _GEN_47;
      end else if (_T_220) begin
        cpr_status_IM_7 <= io_wport_bits_data[15];
      end else begin
        cpr_status_IM_7 <= _GEN_47;
      end
    end else begin
      cpr_status_IM_7 <= _GEN_47;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_UM <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_UM <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_UM <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_UM <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_UM <= _GEN_51;
      end else if (_T_206) begin
        cpr_status_UM <= _GEN_51;
      end else if (_T_211) begin
        cpr_status_UM <= _GEN_51;
      end else if (_T_212) begin
        cpr_status_UM <= _GEN_51;
      end else if (_T_213) begin
        cpr_status_UM <= _GEN_51;
      end else if (_T_219) begin
        cpr_status_UM <= _GEN_51;
      end else if (_T_220) begin
        cpr_status_UM <= io_wport_bits_data[4];
      end else begin
        cpr_status_UM <= _GEN_51;
      end
    end else begin
      cpr_status_UM <= _GEN_51;
    end
    if (io_ex_flush_valid) begin
      if (_T_328) begin
        if (_T_167) begin
          if (_T_168) begin
            if (reset) begin
              cpr_status_ERL <= 1'h0;
            end
          end else if (_T_174) begin
            if (reset) begin
              cpr_status_ERL <= 1'h0;
            end
          end else if (_T_184) begin
            if (reset) begin
              cpr_status_ERL <= 1'h0;
            end
          end else if (_T_194) begin
            if (reset) begin
              cpr_status_ERL <= 1'h0;
            end
          end else if (_T_200) begin
            cpr_status_ERL <= _GEN_53;
          end else if (_T_206) begin
            cpr_status_ERL <= _GEN_53;
          end else if (_T_211) begin
            cpr_status_ERL <= _GEN_53;
          end else if (_T_212) begin
            cpr_status_ERL <= _GEN_53;
          end else if (_T_213) begin
            cpr_status_ERL <= _GEN_53;
          end else if (_T_219) begin
            cpr_status_ERL <= _GEN_53;
          end else if (_T_220) begin
            cpr_status_ERL <= io_wport_bits_data[2];
          end else begin
            cpr_status_ERL <= _GEN_53;
          end
        end else begin
          cpr_status_ERL <= _GEN_53;
        end
      end else if (_T_365) begin
        cpr_status_ERL <= 1'h0;
      end else if (_T_167) begin
        if (_T_168) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_174) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_184) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_194) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_200) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_206) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_211) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_212) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_213) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_219) begin
          cpr_status_ERL <= _GEN_53;
        end else if (_T_220) begin
          cpr_status_ERL <= io_wport_bits_data[2];
        end else begin
          cpr_status_ERL <= _GEN_53;
        end
      end else begin
        cpr_status_ERL <= _GEN_53;
      end
    end else if (_T_167) begin
      if (_T_168) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_174) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_184) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_194) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_200) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_206) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_211) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_212) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_213) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_219) begin
        cpr_status_ERL <= _GEN_53;
      end else if (_T_220) begin
        cpr_status_ERL <= io_wport_bits_data[2];
      end else begin
        cpr_status_ERL <= _GEN_53;
      end
    end else begin
      cpr_status_ERL <= _GEN_53;
    end
    if (io_ex_flush_valid) begin
      if (_T_328) begin
        cpr_status_EXL <= _T_350;
      end else if (_T_167) begin
        if (_T_168) begin
          if (reset) begin
            cpr_status_EXL <= 1'h0;
          end
        end else if (_T_174) begin
          if (reset) begin
            cpr_status_EXL <= 1'h0;
          end
        end else if (_T_184) begin
          if (reset) begin
            cpr_status_EXL <= 1'h0;
          end
        end else if (_T_194) begin
          if (reset) begin
            cpr_status_EXL <= 1'h0;
          end
        end else if (_T_200) begin
          cpr_status_EXL <= _GEN_54;
        end else if (_T_206) begin
          cpr_status_EXL <= _GEN_54;
        end else if (_T_211) begin
          cpr_status_EXL <= _GEN_54;
        end else if (_T_212) begin
          cpr_status_EXL <= _GEN_54;
        end else if (_T_213) begin
          cpr_status_EXL <= _GEN_54;
        end else if (_T_219) begin
          cpr_status_EXL <= _GEN_54;
        end else if (_T_220) begin
          cpr_status_EXL <= io_wport_bits_data[1];
        end else begin
          cpr_status_EXL <= _GEN_54;
        end
      end else begin
        cpr_status_EXL <= _GEN_54;
      end
    end else if (_T_167) begin
      if (_T_168) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_174) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_184) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_194) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_200) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_206) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_211) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_212) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_213) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_219) begin
        cpr_status_EXL <= _GEN_54;
      end else if (_T_220) begin
        cpr_status_EXL <= io_wport_bits_data[1];
      end else begin
        cpr_status_EXL <= _GEN_54;
      end
    end else begin
      cpr_status_EXL <= _GEN_54;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_status_IE <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_status_IE <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_status_IE <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_status_IE <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_status_IE <= _GEN_55;
      end else if (_T_206) begin
        cpr_status_IE <= _GEN_55;
      end else if (_T_211) begin
        cpr_status_IE <= _GEN_55;
      end else if (_T_212) begin
        cpr_status_IE <= _GEN_55;
      end else if (_T_213) begin
        cpr_status_IE <= _GEN_55;
      end else if (_T_219) begin
        cpr_status_IE <= _GEN_55;
      end else if (_T_220) begin
        cpr_status_IE <= io_wport_bits_data[0];
      end else begin
        cpr_status_IE <= _GEN_55;
      end
    end else begin
      cpr_status_IE <= _GEN_55;
    end
    if (io_ex_flush_valid) begin
      if (_T_350) begin
        if (_T_329) begin
          if (is_intr_ex) begin
            cpr_cause_BD <= io_ehu_wb_is_br;
          end else begin
            cpr_cause_BD <= io_ehu_wb_is_ds;
          end
        end else if (reset) begin
          cpr_cause_BD <= 1'h0;
        end
      end else if (reset) begin
        cpr_cause_BD <= 1'h0;
      end
    end else if (reset) begin
      cpr_cause_BD <= 1'h0;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_cause_IV <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_cause_IV <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_cause_IV <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_cause_IV <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_206) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_211) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_212) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_213) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_219) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_220) begin
        cpr_cause_IV <= _GEN_69;
      end else if (_T_251) begin
        cpr_cause_IV <= io_wport_bits_data[23];
      end else begin
        cpr_cause_IV <= _GEN_69;
      end
    end else begin
      cpr_cause_IV <= _GEN_69;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_cause_WP <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_cause_WP <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_cause_WP <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_cause_WP <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_206) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_211) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_212) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_213) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_219) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_220) begin
        cpr_cause_WP <= _GEN_68;
      end else if (_T_251) begin
        cpr_cause_WP <= io_wport_bits_data[22];
      end else begin
        cpr_cause_WP <= _GEN_68;
      end
    end else begin
      cpr_cause_WP <= _GEN_68;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_cause_IP_0 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_cause_IP_0 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_cause_IP_0 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_cause_IP_0 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_206) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_211) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_212) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_213) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_219) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_220) begin
        cpr_cause_IP_0 <= _GEN_59;
      end else if (_T_251) begin
        cpr_cause_IP_0 <= io_wport_bits_data[8];
      end else begin
        cpr_cause_IP_0 <= _GEN_59;
      end
    end else begin
      cpr_cause_IP_0 <= _GEN_59;
    end
    if (_T_167) begin
      if (_T_168) begin
        if (reset) begin
          cpr_cause_IP_1 <= 1'h0;
        end
      end else if (_T_174) begin
        if (reset) begin
          cpr_cause_IP_1 <= 1'h0;
        end
      end else if (_T_184) begin
        if (reset) begin
          cpr_cause_IP_1 <= 1'h0;
        end
      end else if (_T_194) begin
        if (reset) begin
          cpr_cause_IP_1 <= 1'h0;
        end
      end else if (_T_200) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_206) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_211) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_212) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_213) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_219) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_220) begin
        cpr_cause_IP_1 <= _GEN_60;
      end else if (_T_251) begin
        cpr_cause_IP_1 <= io_wport_bits_data[9];
      end else begin
        cpr_cause_IP_1 <= _GEN_60;
      end
    end else begin
      cpr_cause_IP_1 <= _GEN_60;
    end
    cpr_cause_IP_7 <= _T_388 | _GEN_490;
    if (io_ex_flush_valid) begin
      if (_T_350) begin
        if (_T_361) begin
          cpr_cause_ExcCode <= 5'h0;
        end else begin
          cpr_cause_ExcCode <= io_ehu_ex_code;
        end
      end else if (reset) begin
        cpr_cause_ExcCode <= 5'h0;
      end
    end else if (reset) begin
      cpr_cause_ExcCode <= 5'h0;
    end
    if (reset) begin
      cpr_epc <= 32'h0;
    end else if (io_ex_flush_valid) begin
      if (_T_350) begin
        if (_T_329) begin
          if (_T_353) begin
            cpr_epc <= io_ehu_wb_pc;
          end else if (_T_355) begin
            cpr_epc <= io_ehu_wb_npc;
          end else if (io_ehu_wb_is_ds) begin
            cpr_epc <= _T_357;
          end else begin
            cpr_epc <= io_ehu_wb_pc;
          end
        end else if (_T_167) begin
          if (!(_T_168)) begin
            if (!(_T_174)) begin
              if (!(_T_184)) begin
                if (!(_T_194)) begin
                  if (!(_T_200)) begin
                    if (!(_T_206)) begin
                      if (!(_T_211)) begin
                        if (!(_T_212)) begin
                          if (!(_T_213)) begin
                            if (!(_T_219)) begin
                              if (!(_T_220)) begin
                                if (!(_T_251)) begin
                                  if (_T_272) begin
                                    cpr_epc <= io_wport_bits_data;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else if (_T_167) begin
        if (!(_T_168)) begin
          if (!(_T_174)) begin
            if (!(_T_184)) begin
              if (!(_T_194)) begin
                if (!(_T_200)) begin
                  if (!(_T_206)) begin
                    if (!(_T_211)) begin
                      if (!(_T_212)) begin
                        if (!(_T_213)) begin
                          if (!(_T_219)) begin
                            if (!(_T_220)) begin
                              if (!(_T_251)) begin
                                if (_T_272) begin
                                  cpr_epc <= io_wport_bits_data;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else if (_T_167) begin
      if (!(_T_168)) begin
        if (!(_T_174)) begin
          if (!(_T_184)) begin
            if (!(_T_194)) begin
              if (!(_T_200)) begin
                if (!(_T_206)) begin
                  if (!(_T_211)) begin
                    if (!(_T_212)) begin
                      if (!(_T_213)) begin
                        if (!(_T_219)) begin
                          if (!(_T_220)) begin
                            if (!(_T_251)) begin
                              if (_T_272) begin
                                cpr_epc <= io_wport_bits_data;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cpr_ebase <= 32'h0;
    end else if (_T_167) begin
      if (!(_T_168)) begin
        if (!(_T_174)) begin
          if (!(_T_184)) begin
            if (!(_T_194)) begin
              if (!(_T_200)) begin
                if (!(_T_206)) begin
                  if (!(_T_211)) begin
                    if (!(_T_212)) begin
                      if (!(_T_213)) begin
                        if (!(_T_219)) begin
                          if (!(_T_220)) begin
                            if (!(_T_251)) begin
                              if (!(_T_272)) begin
                                if (!(_T_273)) begin
                                  if (_T_274) begin
                                    cpr_ebase <= io_wport_bits_data;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_iaddr_req_ready,
  input         io_iaddr_req_valid,
  input  [31:0] io_iaddr_req_bits_vaddr,
  input         io_iaddr_resp_ready,
  output        io_iaddr_resp_valid,
  output [31:0] io_iaddr_resp_bits_paddr,
  output        io_iaddr_resp_bits_is_cached,
  output [4:0]  io_iaddr_resp_bits_ex_et,
  output [4:0]  io_iaddr_resp_bits_ex_code,
  output [31:0] io_iaddr_resp_bits_ex_addr,
  output [7:0]  io_iaddr_resp_bits_ex_asid,
  output        io_daddr_req_ready,
  input         io_daddr_req_valid,
  input         io_daddr_req_bits_func,
  input  [31:0] io_daddr_req_bits_vaddr,
  input  [1:0]  io_daddr_req_bits_len,
  input         io_daddr_req_bits_is_aligned,
  output [31:0] io_daddr_resp_bits_paddr,
  output [4:0]  io_daddr_resp_bits_ex_et,
  output [4:0]  io_daddr_resp_bits_ex_code,
  output [31:0] io_daddr_resp_bits_ex_addr,
  output [7:0]  io_daddr_resp_bits_ex_asid,
  input  [4:0]  io_rport_index,
  output [15:0] io_rport_entry_pagemask,
  output [18:0] io_rport_entry_vpn,
  output        io_rport_entry_g,
  output [7:0]  io_rport_entry_asid,
  output [23:0] io_rport_entry_p0_pfn,
  output [2:0]  io_rport_entry_p0_c,
  output        io_rport_entry_p0_d,
  output        io_rport_entry_p0_v,
  output [23:0] io_rport_entry_p1_pfn,
  output [2:0]  io_rport_entry_p1_c,
  output        io_rport_entry_p1_d,
  output        io_rport_entry_p1_v,
  input         io_wport_valid,
  input  [4:0]  io_wport_bits_index,
  input  [15:0] io_wport_bits_entry_pagemask,
  input  [18:0] io_wport_bits_entry_vpn,
  input         io_wport_bits_entry_g,
  input  [7:0]  io_wport_bits_entry_asid,
  input  [23:0] io_wport_bits_entry_p0_pfn,
  input  [2:0]  io_wport_bits_entry_p0_c,
  input         io_wport_bits_entry_p0_d,
  input         io_wport_bits_entry_p0_v,
  input  [23:0] io_wport_bits_entry_p1_pfn,
  input  [2:0]  io_wport_bits_entry_p1_c,
  input         io_wport_bits_entry_p1_d,
  input         io_wport_bits_entry_p1_v,
  input  [18:0] io_pport_entry_hi_vpn,
  input  [7:0]  io_pport_entry_hi_asid,
  output        io_pport_index_p,
  output [4:0]  io_pport_index_index,
  input         io_status_ERL,
  input         io_br_flush_valid,
  input         io_ex_flush_valid
);
  reg [15:0] tlb_entries_pagemask [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_0;
  wire [15:0] tlb_entries_pagemask__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_5_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_6_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_7_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_8_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_9_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_10_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_11_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_12_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_13_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_14_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_15_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_16_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_17_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_18_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_19_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_20_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_21_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_22_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_23_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_24_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_25_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_26_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_27_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_28_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_29_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_30_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_31_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_32_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_33_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_34_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_35_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_36_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1546_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1547_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1548_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1549_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1550_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1551_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1552_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1553_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1554_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1555_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1556_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1557_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1558_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1559_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1560_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1561_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1562_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1563_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1564_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1565_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1566_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1567_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1568_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1569_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1570_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1571_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1572_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1573_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1574_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1575_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1576_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask__T_1577_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [15:0] tlb_entries_pagemask_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_pagemask_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_pagemask_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg [18:0] tlb_entries_vpn [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_1;
  wire [18:0] tlb_entries_vpn__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_5_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_6_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_7_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_8_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_9_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_10_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_11_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_12_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_13_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_14_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_15_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_16_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_17_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_18_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_19_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_20_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_21_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_22_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_23_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_24_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_25_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_26_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_27_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_28_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_29_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_30_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_31_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_32_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_33_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_34_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_35_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_36_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1546_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1547_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1548_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1549_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1550_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1551_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1552_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1553_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1554_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1555_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1556_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1557_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1558_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1559_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1560_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1561_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1562_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1563_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1564_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1565_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1566_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1567_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1568_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1569_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1570_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1571_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1572_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1573_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1574_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1575_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1576_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn__T_1577_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [18:0] tlb_entries_vpn_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_vpn_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_vpn_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg  tlb_entries_g [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_2;
  wire  tlb_entries_g__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_5_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_6_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_7_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_8_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_9_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_10_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_11_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_12_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_13_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_14_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_15_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_16_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_17_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_18_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_19_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_20_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_21_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_22_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_23_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_24_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_25_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_26_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_27_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_28_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_29_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_30_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_31_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_32_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_33_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_34_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_35_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_36_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1546_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1547_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1548_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1549_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1550_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1551_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1552_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1553_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1554_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1555_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1556_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1557_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1558_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1559_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1560_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1561_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1562_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1563_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1564_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1565_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1566_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1567_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1568_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1569_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1570_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1571_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1572_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1573_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1574_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1575_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1576_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g__T_1577_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_g_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_g_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg [7:0] tlb_entries_asid [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_3;
  wire [7:0] tlb_entries_asid__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_5_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_6_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_7_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_8_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_9_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_10_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_11_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_12_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_13_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_14_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_15_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_16_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_17_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_18_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_19_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_20_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_21_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_22_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_23_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_24_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_25_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_26_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_27_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_28_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_29_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_30_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_31_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_32_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_33_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_34_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_35_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_36_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1546_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1547_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1548_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1549_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1550_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1551_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1552_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1553_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1554_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1555_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1556_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1557_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1558_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1559_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1560_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1561_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1562_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1563_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1564_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1565_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1566_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1567_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1568_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1569_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1570_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1571_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1572_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1573_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1574_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1575_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1576_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid__T_1577_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [7:0] tlb_entries_asid_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_asid_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_asid_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg [23:0] tlb_entries_p0_pfn [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_4;
  wire [23:0] tlb_entries_p0_pfn__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_5_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_6_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_7_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_8_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_9_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_10_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_11_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_12_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_13_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_14_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_15_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_16_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_17_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_18_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_19_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_20_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_21_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_22_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_23_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_24_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_25_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_26_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_27_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_28_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_29_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_30_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_31_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_32_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_33_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_34_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_35_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_36_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1546_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1547_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1548_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1549_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1550_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1551_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1552_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1553_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1554_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1555_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1556_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1557_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1558_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1559_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1560_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1561_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1562_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1563_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1564_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1565_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1566_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1567_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1568_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1569_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1570_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1571_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1572_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1573_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1574_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1575_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1576_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn__T_1577_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p0_pfn_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_pfn_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_pfn_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg [2:0] tlb_entries_p0_c [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_5;
  wire [2:0] tlb_entries_p0_c__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_5_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_6_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_7_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_8_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_9_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_10_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_11_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_12_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_13_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_14_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_15_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_16_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_17_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_18_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_19_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_20_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_21_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_22_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_23_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_24_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_25_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_26_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_27_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_28_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_29_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_30_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_31_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_32_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_33_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_34_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_35_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_36_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1546_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1547_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1548_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1549_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1550_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1551_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1552_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1553_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1554_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1555_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1556_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1557_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1558_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1559_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1560_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1561_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1562_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1563_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1564_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1565_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1566_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1567_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1568_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1569_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1570_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1571_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1572_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1573_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1574_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1575_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1576_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c__T_1577_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p0_c_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_c_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_c_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg  tlb_entries_p0_d [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_6;
  wire  tlb_entries_p0_d__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_5_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_6_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_7_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_8_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_9_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_10_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_11_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_12_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_13_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_14_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_15_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_16_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_17_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_18_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_19_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_20_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_21_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_22_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_23_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_24_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_25_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_26_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_27_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_28_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_29_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_30_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_31_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_32_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_33_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_34_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_35_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_36_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1546_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1547_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1548_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1549_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1550_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1551_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1552_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1553_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1554_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1555_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1556_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1557_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1558_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1559_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1560_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1561_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1562_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1563_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1564_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1565_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1566_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1567_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1568_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1569_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1570_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1571_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1572_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1573_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1574_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1575_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1576_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d__T_1577_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_d_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_d_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg  tlb_entries_p0_v [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_7;
  wire  tlb_entries_p0_v__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_5_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_6_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_7_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_8_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_9_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_10_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_11_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_12_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_13_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_14_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_15_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_16_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_17_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_18_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_19_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_20_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_21_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_22_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_23_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_24_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_25_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_26_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_27_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_28_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_29_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_30_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_31_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_32_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_33_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_34_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_35_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_36_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1546_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1547_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1548_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1549_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1550_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1551_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1552_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1553_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1554_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1555_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1556_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1557_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1558_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1559_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1560_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1561_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1562_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1563_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1564_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1565_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1566_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1567_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1568_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1569_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1570_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1571_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1572_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1573_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1574_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1575_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1576_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v__T_1577_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p0_v_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p0_v_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg [23:0] tlb_entries_p1_pfn [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_8;
  wire [23:0] tlb_entries_p1_pfn__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_5_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_6_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_7_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_8_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_9_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_10_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_11_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_12_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_13_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_14_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_15_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_16_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_17_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_18_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_19_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_20_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_21_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_22_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_23_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_24_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_25_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_26_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_27_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_28_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_29_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_30_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_31_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_32_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_33_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_34_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_35_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_36_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1546_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1547_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1548_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1549_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1550_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1551_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1552_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1553_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1554_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1555_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1556_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1557_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1558_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1559_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1560_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1561_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1562_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1563_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1564_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1565_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1566_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1567_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1568_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1569_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1570_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1571_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1572_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1573_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1574_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1575_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1576_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn__T_1577_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [23:0] tlb_entries_p1_pfn_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_pfn_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_pfn_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg [2:0] tlb_entries_p1_c [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_9;
  wire [2:0] tlb_entries_p1_c__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_5_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_6_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_7_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_8_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_9_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_10_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_11_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_12_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_13_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_14_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_15_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_16_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_17_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_18_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_19_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_20_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_21_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_22_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_23_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_24_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_25_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_26_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_27_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_28_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_29_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_30_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_31_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_32_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_33_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_34_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_35_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_36_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1546_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1547_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1548_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1549_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1550_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1551_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1552_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1553_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1554_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1555_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1556_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1557_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1558_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1559_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1560_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1561_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1562_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1563_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1564_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1565_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1566_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1567_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1568_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1569_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1570_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1571_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1572_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1573_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1574_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1575_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1576_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c__T_1577_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire [2:0] tlb_entries_p1_c_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_c_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_c_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg  tlb_entries_p1_d [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_10;
  wire  tlb_entries_p1_d__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_5_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_6_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_7_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_8_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_9_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_10_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_11_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_12_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_13_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_14_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_15_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_16_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_17_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_18_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_19_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_20_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_21_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_22_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_23_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_24_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_25_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_26_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_27_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_28_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_29_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_30_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_31_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_32_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_33_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_34_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_35_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_36_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1546_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1547_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1548_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1549_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1550_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1551_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1552_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1553_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1554_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1555_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1556_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1557_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1558_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1559_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1560_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1561_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1562_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1563_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1564_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1565_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1566_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1567_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1568_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1569_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1570_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1571_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1572_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1573_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1574_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1575_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1576_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d__T_1577_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_d_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_d_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  reg  tlb_entries_p1_v [0:31]; // @[tlb.scala 45:24]
  reg [31:0] _RAND_11;
  wire  tlb_entries_p1_v__T_5_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_5_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_6_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_6_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_7_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_7_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_8_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_8_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_9_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_9_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_10_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_10_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_11_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_11_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_12_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_12_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_13_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_13_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_14_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_14_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_15_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_15_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_16_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_16_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_17_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_17_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_18_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_18_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_19_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_19_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_20_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_20_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_21_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_21_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_22_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_22_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_23_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_23_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_24_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_24_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_25_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_25_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_26_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_26_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_27_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_27_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_28_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_28_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_29_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_29_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_30_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_30_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_31_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_31_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_32_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_32_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_33_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_33_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_34_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_34_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_35_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_35_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_36_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_36_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1546_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1546_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1547_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1547_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1548_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1548_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1549_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1549_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1550_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1550_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1551_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1551_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1552_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1552_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1553_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1553_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1554_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1554_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1555_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1555_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1556_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1556_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1557_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1557_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1558_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1558_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1559_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1559_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1560_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1560_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1561_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1561_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1562_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1562_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1563_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1563_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1564_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1564_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1565_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1565_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1566_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1566_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1567_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1567_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1568_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1568_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1569_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1569_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1570_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1570_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1571_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1571_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1572_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1572_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1573_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1573_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1574_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1574_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1575_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1575_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1576_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1576_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v__T_1577_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v__T_1577_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_0_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_0_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_1_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_1_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_2_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_2_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_3_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_3_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_4_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_4_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_5_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_5_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_6_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_6_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_7_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_7_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_8_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_8_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_9_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_9_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_10_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_10_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_11_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_11_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_12_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_12_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_13_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_13_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_14_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_14_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_15_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_15_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_16_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_16_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_17_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_17_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_18_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_18_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_19_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_19_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_20_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_20_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_21_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_21_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_22_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_22_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_23_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_23_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_24_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_24_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_25_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_25_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_26_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_26_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_27_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_27_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_28_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_28_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_29_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_29_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_30_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_30_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_31_r_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_31_r_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_0_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_0_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_0_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_1_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_1_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_1_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_2_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_2_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_2_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_3_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_3_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_3_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_4_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_4_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_4_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_5_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_5_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_5_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_6_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_6_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_6_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_7_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_7_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_7_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_8_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_8_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_8_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_9_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_9_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_9_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_10_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_10_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_10_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_11_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_11_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_11_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_12_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_12_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_12_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_13_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_13_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_13_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_14_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_14_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_14_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_15_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_15_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_15_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_16_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_16_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_16_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_17_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_17_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_17_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_18_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_18_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_18_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_19_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_19_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_19_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_20_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_20_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_20_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_21_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_21_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_21_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_22_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_22_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_22_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_23_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_23_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_23_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_24_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_24_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_24_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_25_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_25_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_25_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_26_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_26_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_26_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_27_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_27_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_27_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_28_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_28_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_28_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_29_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_29_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_29_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_30_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_30_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_30_w_en; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
  wire [4:0] tlb_entries_p1_v_tlb_entry_ports_31_w_addr; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_31_w_mask; // @[tlb.scala 45:24]
  wire  tlb_entries_p1_v_tlb_entry_ports_31_w_en; // @[tlb.scala 45:24]
  wire  _T = io_br_flush_valid | io_ex_flush_valid; // @[tlb.scala 185:60]
  wire  _T_1 = io_iaddr_req_ready & io_iaddr_req_valid; // @[Decoupled.scala 40:37]
  reg [31:0] _T_3_vaddr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg [1:0] _T_3_len; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg  _T_3_is_aligned; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  wire  _GEN_0 = _T_1 | _T_3_is_aligned; // @[Reg.scala 28:19]
  reg  _T_4; // @[tlb.scala 146:31]
  reg [31:0] _RAND_15;
  wire [31:0] _T_38 = {{16'd0}, tlb_entries_pagemask__T_5_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_39 = ~_T_38; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1228 = {{13'd0}, tlb_entries_vpn__T_5_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_40 = _GEN_1228 & _T_39; // @[tlb.scala 50:19]
  wire [31:0] _GEN_1229 = {{13'd0}, _T_3_vaddr[31:13]}; // @[tlb.scala 50:37]
  wire [31:0] _T_42 = _GEN_1229 & _T_39; // @[tlb.scala 50:37]
  wire  _T_43 = _T_40 == _T_42; // @[tlb.scala 50:28]
  wire  _T_44 = tlb_entries_asid__T_5_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_45 = tlb_entries_g__T_5_data | _T_44; // @[tlb.scala 51:17]
  wire  _T_46 = _T_43 & _T_45; // @[tlb.scala 50:46]
  wire [31:0] _T_48 = {{16'd0}, tlb_entries_pagemask__T_6_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_49 = ~_T_48; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1230 = {{13'd0}, tlb_entries_vpn__T_6_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_50 = _GEN_1230 & _T_49; // @[tlb.scala 50:19]
  wire [31:0] _T_52 = _GEN_1229 & _T_49; // @[tlb.scala 50:37]
  wire  _T_53 = _T_50 == _T_52; // @[tlb.scala 50:28]
  wire  _T_54 = tlb_entries_asid__T_6_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_55 = tlb_entries_g__T_6_data | _T_54; // @[tlb.scala 51:17]
  wire  _T_56 = _T_53 & _T_55; // @[tlb.scala 50:46]
  wire [31:0] _T_58 = {{16'd0}, tlb_entries_pagemask__T_7_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_59 = ~_T_58; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1232 = {{13'd0}, tlb_entries_vpn__T_7_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_60 = _GEN_1232 & _T_59; // @[tlb.scala 50:19]
  wire [31:0] _T_62 = _GEN_1229 & _T_59; // @[tlb.scala 50:37]
  wire  _T_63 = _T_60 == _T_62; // @[tlb.scala 50:28]
  wire  _T_64 = tlb_entries_asid__T_7_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_65 = tlb_entries_g__T_7_data | _T_64; // @[tlb.scala 51:17]
  wire  _T_66 = _T_63 & _T_65; // @[tlb.scala 50:46]
  wire [31:0] _T_68 = {{16'd0}, tlb_entries_pagemask__T_8_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_69 = ~_T_68; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1234 = {{13'd0}, tlb_entries_vpn__T_8_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_70 = _GEN_1234 & _T_69; // @[tlb.scala 50:19]
  wire [31:0] _T_72 = _GEN_1229 & _T_69; // @[tlb.scala 50:37]
  wire  _T_73 = _T_70 == _T_72; // @[tlb.scala 50:28]
  wire  _T_74 = tlb_entries_asid__T_8_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_75 = tlb_entries_g__T_8_data | _T_74; // @[tlb.scala 51:17]
  wire  _T_76 = _T_73 & _T_75; // @[tlb.scala 50:46]
  wire [31:0] _T_78 = {{16'd0}, tlb_entries_pagemask__T_9_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_79 = ~_T_78; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1236 = {{13'd0}, tlb_entries_vpn__T_9_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_80 = _GEN_1236 & _T_79; // @[tlb.scala 50:19]
  wire [31:0] _T_82 = _GEN_1229 & _T_79; // @[tlb.scala 50:37]
  wire  _T_83 = _T_80 == _T_82; // @[tlb.scala 50:28]
  wire  _T_84 = tlb_entries_asid__T_9_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_85 = tlb_entries_g__T_9_data | _T_84; // @[tlb.scala 51:17]
  wire  _T_86 = _T_83 & _T_85; // @[tlb.scala 50:46]
  wire [31:0] _T_88 = {{16'd0}, tlb_entries_pagemask__T_10_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_89 = ~_T_88; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1238 = {{13'd0}, tlb_entries_vpn__T_10_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_90 = _GEN_1238 & _T_89; // @[tlb.scala 50:19]
  wire [31:0] _T_92 = _GEN_1229 & _T_89; // @[tlb.scala 50:37]
  wire  _T_93 = _T_90 == _T_92; // @[tlb.scala 50:28]
  wire  _T_94 = tlb_entries_asid__T_10_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_95 = tlb_entries_g__T_10_data | _T_94; // @[tlb.scala 51:17]
  wire  _T_96 = _T_93 & _T_95; // @[tlb.scala 50:46]
  wire [31:0] _T_98 = {{16'd0}, tlb_entries_pagemask__T_11_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_99 = ~_T_98; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1240 = {{13'd0}, tlb_entries_vpn__T_11_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_100 = _GEN_1240 & _T_99; // @[tlb.scala 50:19]
  wire [31:0] _T_102 = _GEN_1229 & _T_99; // @[tlb.scala 50:37]
  wire  _T_103 = _T_100 == _T_102; // @[tlb.scala 50:28]
  wire  _T_104 = tlb_entries_asid__T_11_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_105 = tlb_entries_g__T_11_data | _T_104; // @[tlb.scala 51:17]
  wire  _T_106 = _T_103 & _T_105; // @[tlb.scala 50:46]
  wire [31:0] _T_108 = {{16'd0}, tlb_entries_pagemask__T_12_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_109 = ~_T_108; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1242 = {{13'd0}, tlb_entries_vpn__T_12_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_110 = _GEN_1242 & _T_109; // @[tlb.scala 50:19]
  wire [31:0] _T_112 = _GEN_1229 & _T_109; // @[tlb.scala 50:37]
  wire  _T_113 = _T_110 == _T_112; // @[tlb.scala 50:28]
  wire  _T_114 = tlb_entries_asid__T_12_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_115 = tlb_entries_g__T_12_data | _T_114; // @[tlb.scala 51:17]
  wire  _T_116 = _T_113 & _T_115; // @[tlb.scala 50:46]
  wire [31:0] _T_118 = {{16'd0}, tlb_entries_pagemask__T_13_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_119 = ~_T_118; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1244 = {{13'd0}, tlb_entries_vpn__T_13_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_120 = _GEN_1244 & _T_119; // @[tlb.scala 50:19]
  wire [31:0] _T_122 = _GEN_1229 & _T_119; // @[tlb.scala 50:37]
  wire  _T_123 = _T_120 == _T_122; // @[tlb.scala 50:28]
  wire  _T_124 = tlb_entries_asid__T_13_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_125 = tlb_entries_g__T_13_data | _T_124; // @[tlb.scala 51:17]
  wire  _T_126 = _T_123 & _T_125; // @[tlb.scala 50:46]
  wire [31:0] _T_128 = {{16'd0}, tlb_entries_pagemask__T_14_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_129 = ~_T_128; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1246 = {{13'd0}, tlb_entries_vpn__T_14_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_130 = _GEN_1246 & _T_129; // @[tlb.scala 50:19]
  wire [31:0] _T_132 = _GEN_1229 & _T_129; // @[tlb.scala 50:37]
  wire  _T_133 = _T_130 == _T_132; // @[tlb.scala 50:28]
  wire  _T_134 = tlb_entries_asid__T_14_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_135 = tlb_entries_g__T_14_data | _T_134; // @[tlb.scala 51:17]
  wire  _T_136 = _T_133 & _T_135; // @[tlb.scala 50:46]
  wire [31:0] _T_138 = {{16'd0}, tlb_entries_pagemask__T_15_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_139 = ~_T_138; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1248 = {{13'd0}, tlb_entries_vpn__T_15_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_140 = _GEN_1248 & _T_139; // @[tlb.scala 50:19]
  wire [31:0] _T_142 = _GEN_1229 & _T_139; // @[tlb.scala 50:37]
  wire  _T_143 = _T_140 == _T_142; // @[tlb.scala 50:28]
  wire  _T_144 = tlb_entries_asid__T_15_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_145 = tlb_entries_g__T_15_data | _T_144; // @[tlb.scala 51:17]
  wire  _T_146 = _T_143 & _T_145; // @[tlb.scala 50:46]
  wire [31:0] _T_148 = {{16'd0}, tlb_entries_pagemask__T_16_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_149 = ~_T_148; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1250 = {{13'd0}, tlb_entries_vpn__T_16_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_150 = _GEN_1250 & _T_149; // @[tlb.scala 50:19]
  wire [31:0] _T_152 = _GEN_1229 & _T_149; // @[tlb.scala 50:37]
  wire  _T_153 = _T_150 == _T_152; // @[tlb.scala 50:28]
  wire  _T_154 = tlb_entries_asid__T_16_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_155 = tlb_entries_g__T_16_data | _T_154; // @[tlb.scala 51:17]
  wire  _T_156 = _T_153 & _T_155; // @[tlb.scala 50:46]
  wire [31:0] _T_158 = {{16'd0}, tlb_entries_pagemask__T_17_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_159 = ~_T_158; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1252 = {{13'd0}, tlb_entries_vpn__T_17_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_160 = _GEN_1252 & _T_159; // @[tlb.scala 50:19]
  wire [31:0] _T_162 = _GEN_1229 & _T_159; // @[tlb.scala 50:37]
  wire  _T_163 = _T_160 == _T_162; // @[tlb.scala 50:28]
  wire  _T_164 = tlb_entries_asid__T_17_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_165 = tlb_entries_g__T_17_data | _T_164; // @[tlb.scala 51:17]
  wire  _T_166 = _T_163 & _T_165; // @[tlb.scala 50:46]
  wire [31:0] _T_168 = {{16'd0}, tlb_entries_pagemask__T_18_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_169 = ~_T_168; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1254 = {{13'd0}, tlb_entries_vpn__T_18_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_170 = _GEN_1254 & _T_169; // @[tlb.scala 50:19]
  wire [31:0] _T_172 = _GEN_1229 & _T_169; // @[tlb.scala 50:37]
  wire  _T_173 = _T_170 == _T_172; // @[tlb.scala 50:28]
  wire  _T_174 = tlb_entries_asid__T_18_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_175 = tlb_entries_g__T_18_data | _T_174; // @[tlb.scala 51:17]
  wire  _T_176 = _T_173 & _T_175; // @[tlb.scala 50:46]
  wire [31:0] _T_178 = {{16'd0}, tlb_entries_pagemask__T_19_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_179 = ~_T_178; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1256 = {{13'd0}, tlb_entries_vpn__T_19_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_180 = _GEN_1256 & _T_179; // @[tlb.scala 50:19]
  wire [31:0] _T_182 = _GEN_1229 & _T_179; // @[tlb.scala 50:37]
  wire  _T_183 = _T_180 == _T_182; // @[tlb.scala 50:28]
  wire  _T_184 = tlb_entries_asid__T_19_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_185 = tlb_entries_g__T_19_data | _T_184; // @[tlb.scala 51:17]
  wire  _T_186 = _T_183 & _T_185; // @[tlb.scala 50:46]
  wire [31:0] _T_188 = {{16'd0}, tlb_entries_pagemask__T_20_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_189 = ~_T_188; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1258 = {{13'd0}, tlb_entries_vpn__T_20_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_190 = _GEN_1258 & _T_189; // @[tlb.scala 50:19]
  wire [31:0] _T_192 = _GEN_1229 & _T_189; // @[tlb.scala 50:37]
  wire  _T_193 = _T_190 == _T_192; // @[tlb.scala 50:28]
  wire  _T_194 = tlb_entries_asid__T_20_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_195 = tlb_entries_g__T_20_data | _T_194; // @[tlb.scala 51:17]
  wire  _T_196 = _T_193 & _T_195; // @[tlb.scala 50:46]
  wire [31:0] _T_198 = {{16'd0}, tlb_entries_pagemask__T_21_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_199 = ~_T_198; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1260 = {{13'd0}, tlb_entries_vpn__T_21_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_200 = _GEN_1260 & _T_199; // @[tlb.scala 50:19]
  wire [31:0] _T_202 = _GEN_1229 & _T_199; // @[tlb.scala 50:37]
  wire  _T_203 = _T_200 == _T_202; // @[tlb.scala 50:28]
  wire  _T_204 = tlb_entries_asid__T_21_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_205 = tlb_entries_g__T_21_data | _T_204; // @[tlb.scala 51:17]
  wire  _T_206 = _T_203 & _T_205; // @[tlb.scala 50:46]
  wire [31:0] _T_208 = {{16'd0}, tlb_entries_pagemask__T_22_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_209 = ~_T_208; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1262 = {{13'd0}, tlb_entries_vpn__T_22_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_210 = _GEN_1262 & _T_209; // @[tlb.scala 50:19]
  wire [31:0] _T_212 = _GEN_1229 & _T_209; // @[tlb.scala 50:37]
  wire  _T_213 = _T_210 == _T_212; // @[tlb.scala 50:28]
  wire  _T_214 = tlb_entries_asid__T_22_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_215 = tlb_entries_g__T_22_data | _T_214; // @[tlb.scala 51:17]
  wire  _T_216 = _T_213 & _T_215; // @[tlb.scala 50:46]
  wire [31:0] _T_218 = {{16'd0}, tlb_entries_pagemask__T_23_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_219 = ~_T_218; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1264 = {{13'd0}, tlb_entries_vpn__T_23_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_220 = _GEN_1264 & _T_219; // @[tlb.scala 50:19]
  wire [31:0] _T_222 = _GEN_1229 & _T_219; // @[tlb.scala 50:37]
  wire  _T_223 = _T_220 == _T_222; // @[tlb.scala 50:28]
  wire  _T_224 = tlb_entries_asid__T_23_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_225 = tlb_entries_g__T_23_data | _T_224; // @[tlb.scala 51:17]
  wire  _T_226 = _T_223 & _T_225; // @[tlb.scala 50:46]
  wire [31:0] _T_228 = {{16'd0}, tlb_entries_pagemask__T_24_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_229 = ~_T_228; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1266 = {{13'd0}, tlb_entries_vpn__T_24_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_230 = _GEN_1266 & _T_229; // @[tlb.scala 50:19]
  wire [31:0] _T_232 = _GEN_1229 & _T_229; // @[tlb.scala 50:37]
  wire  _T_233 = _T_230 == _T_232; // @[tlb.scala 50:28]
  wire  _T_234 = tlb_entries_asid__T_24_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_235 = tlb_entries_g__T_24_data | _T_234; // @[tlb.scala 51:17]
  wire  _T_236 = _T_233 & _T_235; // @[tlb.scala 50:46]
  wire [31:0] _T_238 = {{16'd0}, tlb_entries_pagemask__T_25_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_239 = ~_T_238; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1268 = {{13'd0}, tlb_entries_vpn__T_25_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_240 = _GEN_1268 & _T_239; // @[tlb.scala 50:19]
  wire [31:0] _T_242 = _GEN_1229 & _T_239; // @[tlb.scala 50:37]
  wire  _T_243 = _T_240 == _T_242; // @[tlb.scala 50:28]
  wire  _T_244 = tlb_entries_asid__T_25_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_245 = tlb_entries_g__T_25_data | _T_244; // @[tlb.scala 51:17]
  wire  _T_246 = _T_243 & _T_245; // @[tlb.scala 50:46]
  wire [31:0] _T_248 = {{16'd0}, tlb_entries_pagemask__T_26_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_249 = ~_T_248; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1270 = {{13'd0}, tlb_entries_vpn__T_26_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_250 = _GEN_1270 & _T_249; // @[tlb.scala 50:19]
  wire [31:0] _T_252 = _GEN_1229 & _T_249; // @[tlb.scala 50:37]
  wire  _T_253 = _T_250 == _T_252; // @[tlb.scala 50:28]
  wire  _T_254 = tlb_entries_asid__T_26_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_255 = tlb_entries_g__T_26_data | _T_254; // @[tlb.scala 51:17]
  wire  _T_256 = _T_253 & _T_255; // @[tlb.scala 50:46]
  wire [31:0] _T_258 = {{16'd0}, tlb_entries_pagemask__T_27_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_259 = ~_T_258; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1272 = {{13'd0}, tlb_entries_vpn__T_27_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_260 = _GEN_1272 & _T_259; // @[tlb.scala 50:19]
  wire [31:0] _T_262 = _GEN_1229 & _T_259; // @[tlb.scala 50:37]
  wire  _T_263 = _T_260 == _T_262; // @[tlb.scala 50:28]
  wire  _T_264 = tlb_entries_asid__T_27_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_265 = tlb_entries_g__T_27_data | _T_264; // @[tlb.scala 51:17]
  wire  _T_266 = _T_263 & _T_265; // @[tlb.scala 50:46]
  wire [31:0] _T_268 = {{16'd0}, tlb_entries_pagemask__T_28_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_269 = ~_T_268; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1274 = {{13'd0}, tlb_entries_vpn__T_28_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_270 = _GEN_1274 & _T_269; // @[tlb.scala 50:19]
  wire [31:0] _T_272 = _GEN_1229 & _T_269; // @[tlb.scala 50:37]
  wire  _T_273 = _T_270 == _T_272; // @[tlb.scala 50:28]
  wire  _T_274 = tlb_entries_asid__T_28_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_275 = tlb_entries_g__T_28_data | _T_274; // @[tlb.scala 51:17]
  wire  _T_276 = _T_273 & _T_275; // @[tlb.scala 50:46]
  wire [31:0] _T_278 = {{16'd0}, tlb_entries_pagemask__T_29_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_279 = ~_T_278; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1276 = {{13'd0}, tlb_entries_vpn__T_29_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_280 = _GEN_1276 & _T_279; // @[tlb.scala 50:19]
  wire [31:0] _T_282 = _GEN_1229 & _T_279; // @[tlb.scala 50:37]
  wire  _T_283 = _T_280 == _T_282; // @[tlb.scala 50:28]
  wire  _T_284 = tlb_entries_asid__T_29_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_285 = tlb_entries_g__T_29_data | _T_284; // @[tlb.scala 51:17]
  wire  _T_286 = _T_283 & _T_285; // @[tlb.scala 50:46]
  wire [31:0] _T_288 = {{16'd0}, tlb_entries_pagemask__T_30_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_289 = ~_T_288; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1278 = {{13'd0}, tlb_entries_vpn__T_30_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_290 = _GEN_1278 & _T_289; // @[tlb.scala 50:19]
  wire [31:0] _T_292 = _GEN_1229 & _T_289; // @[tlb.scala 50:37]
  wire  _T_293 = _T_290 == _T_292; // @[tlb.scala 50:28]
  wire  _T_294 = tlb_entries_asid__T_30_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_295 = tlb_entries_g__T_30_data | _T_294; // @[tlb.scala 51:17]
  wire  _T_296 = _T_293 & _T_295; // @[tlb.scala 50:46]
  wire [31:0] _T_298 = {{16'd0}, tlb_entries_pagemask__T_31_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_299 = ~_T_298; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1280 = {{13'd0}, tlb_entries_vpn__T_31_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_300 = _GEN_1280 & _T_299; // @[tlb.scala 50:19]
  wire [31:0] _T_302 = _GEN_1229 & _T_299; // @[tlb.scala 50:37]
  wire  _T_303 = _T_300 == _T_302; // @[tlb.scala 50:28]
  wire  _T_304 = tlb_entries_asid__T_31_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_305 = tlb_entries_g__T_31_data | _T_304; // @[tlb.scala 51:17]
  wire  _T_306 = _T_303 & _T_305; // @[tlb.scala 50:46]
  wire [31:0] _T_308 = {{16'd0}, tlb_entries_pagemask__T_32_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_309 = ~_T_308; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1282 = {{13'd0}, tlb_entries_vpn__T_32_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_310 = _GEN_1282 & _T_309; // @[tlb.scala 50:19]
  wire [31:0] _T_312 = _GEN_1229 & _T_309; // @[tlb.scala 50:37]
  wire  _T_313 = _T_310 == _T_312; // @[tlb.scala 50:28]
  wire  _T_314 = tlb_entries_asid__T_32_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_315 = tlb_entries_g__T_32_data | _T_314; // @[tlb.scala 51:17]
  wire  _T_316 = _T_313 & _T_315; // @[tlb.scala 50:46]
  wire [31:0] _T_318 = {{16'd0}, tlb_entries_pagemask__T_33_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_319 = ~_T_318; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1284 = {{13'd0}, tlb_entries_vpn__T_33_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_320 = _GEN_1284 & _T_319; // @[tlb.scala 50:19]
  wire [31:0] _T_322 = _GEN_1229 & _T_319; // @[tlb.scala 50:37]
  wire  _T_323 = _T_320 == _T_322; // @[tlb.scala 50:28]
  wire  _T_324 = tlb_entries_asid__T_33_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_325 = tlb_entries_g__T_33_data | _T_324; // @[tlb.scala 51:17]
  wire  _T_326 = _T_323 & _T_325; // @[tlb.scala 50:46]
  wire [31:0] _T_328 = {{16'd0}, tlb_entries_pagemask__T_34_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_329 = ~_T_328; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1286 = {{13'd0}, tlb_entries_vpn__T_34_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_330 = _GEN_1286 & _T_329; // @[tlb.scala 50:19]
  wire [31:0] _T_332 = _GEN_1229 & _T_329; // @[tlb.scala 50:37]
  wire  _T_333 = _T_330 == _T_332; // @[tlb.scala 50:28]
  wire  _T_334 = tlb_entries_asid__T_34_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_335 = tlb_entries_g__T_34_data | _T_334; // @[tlb.scala 51:17]
  wire  _T_336 = _T_333 & _T_335; // @[tlb.scala 50:46]
  wire [31:0] _T_338 = {{16'd0}, tlb_entries_pagemask__T_35_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_339 = ~_T_338; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1288 = {{13'd0}, tlb_entries_vpn__T_35_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_340 = _GEN_1288 & _T_339; // @[tlb.scala 50:19]
  wire [31:0] _T_342 = _GEN_1229 & _T_339; // @[tlb.scala 50:37]
  wire  _T_343 = _T_340 == _T_342; // @[tlb.scala 50:28]
  wire  _T_344 = tlb_entries_asid__T_35_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_345 = tlb_entries_g__T_35_data | _T_344; // @[tlb.scala 51:17]
  wire  _T_346 = _T_343 & _T_345; // @[tlb.scala 50:46]
  wire [31:0] _T_348 = {{16'd0}, tlb_entries_pagemask__T_36_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_349 = ~_T_348; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1290 = {{13'd0}, tlb_entries_vpn__T_36_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_350 = _GEN_1290 & _T_349; // @[tlb.scala 50:19]
  wire [31:0] _T_352 = _GEN_1229 & _T_349; // @[tlb.scala 50:37]
  wire  _T_353 = _T_350 == _T_352; // @[tlb.scala 50:28]
  wire  _T_354 = tlb_entries_asid__T_36_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_355 = tlb_entries_g__T_36_data | _T_354; // @[tlb.scala 51:17]
  wire  _T_356 = _T_353 & _T_355; // @[tlb.scala 50:46]
  wire [7:0] _T_363 = {_T_286,_T_296,_T_306,_T_316,_T_326,_T_336,_T_346,_T_356}; // @[Cat.scala 29:58]
  wire [15:0] _T_371 = {_T_206,_T_216,_T_226,_T_236,_T_246,_T_256,_T_266,_T_276,_T_363}; // @[Cat.scala 29:58]
  wire [7:0] _T_378 = {_T_126,_T_136,_T_146,_T_156,_T_166,_T_176,_T_186,_T_196}; // @[Cat.scala 29:58]
  wire [31:0] _T_387 = {_T_46,_T_56,_T_66,_T_76,_T_86,_T_96,_T_106,_T_116,_T_378,_T_371}; // @[Cat.scala 29:58]
  wire [31:0] _T_391 = {{16'd0}, _T_387[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_393 = {_T_387[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_395 = _T_393 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_396 = _T_391 | _T_395; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1292 = {{8'd0}, _T_396[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_401 = _GEN_1292 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_403 = {_T_396[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_405 = _T_403 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_406 = _T_401 | _T_405; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1293 = {{4'd0}, _T_406[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_411 = _GEN_1293 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_413 = {_T_406[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_415 = _T_413 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_416 = _T_411 | _T_415; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1294 = {{2'd0}, _T_416[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_421 = _GEN_1294 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_423 = {_T_416[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_425 = _T_423 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_426 = _T_421 | _T_425; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1295 = {{1'd0}, _T_426[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_431 = _GEN_1295 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_433 = {_T_426[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_435 = _T_433 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_436 = _T_431 | _T_435; // @[Bitwise.scala 103:39]
  wire  _T_437 = _T_436 != 32'h0; // @[tlb.scala 83:25]
  wire  _T_438 = ~_T_437; // @[tlb.scala 83:16]
  wire [31:0] _T_442 = _T_38 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_443 = {_T_442, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _GEN_1296 = {{12'd0}, _T_3_vaddr}; // @[tlb.scala 55:24]
  wire [43:0] _T_444 = _GEN_1296 & _T_443; // @[tlb.scala 55:24]
  wire  _T_445 = _T_444 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_446_pfn = _T_445 ? tlb_entries_p1_pfn__T_5_data : tlb_entries_p0_pfn__T_5_data; // @[tlb.scala 56:19]
  wire  _T_446_v = _T_445 ? tlb_entries_p1_v__T_5_data : tlb_entries_p0_v__T_5_data; // @[tlb.scala 56:19]
  wire  _T_451 = ~_T_446_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1297 = {{8'd0}, _T_446_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_456 = _GEN_1297 & _T_39; // @[tlb.scala 68:32]
  wire [43:0] _T_457 = {_T_456, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_462 = _T_443 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_463 = _GEN_1296 & _T_462; // @[tlb.scala 69:27]
  wire [43:0] _T_464 = _T_457 | _T_463; // @[tlb.scala 70:29]
  wire [4:0] _GEN_7 = _T_451 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_9 = _T_451 ? 44'h0 : _T_464; // @[tlb.scala 59:27]
  wire [31:0] _T_468 = _T_48 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_469 = {_T_468, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_470 = _GEN_1296 & _T_469; // @[tlb.scala 55:24]
  wire  _T_471 = _T_470 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_472_pfn = _T_471 ? tlb_entries_p1_pfn__T_6_data : tlb_entries_p0_pfn__T_6_data; // @[tlb.scala 56:19]
  wire  _T_472_v = _T_471 ? tlb_entries_p1_v__T_6_data : tlb_entries_p0_v__T_6_data; // @[tlb.scala 56:19]
  wire  _T_477 = ~_T_472_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1300 = {{8'd0}, _T_472_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_482 = _GEN_1300 & _T_49; // @[tlb.scala 68:32]
  wire [43:0] _T_483 = {_T_482, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_488 = _T_469 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_489 = _GEN_1296 & _T_488; // @[tlb.scala 69:27]
  wire [43:0] _T_490 = _T_483 | _T_489; // @[tlb.scala 70:29]
  wire [4:0] _GEN_13 = _T_477 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_15 = _T_477 ? 44'h0 : _T_490; // @[tlb.scala 59:27]
  wire [31:0] _T_494 = _T_58 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_495 = {_T_494, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_496 = _GEN_1296 & _T_495; // @[tlb.scala 55:24]
  wire  _T_497 = _T_496 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_498_pfn = _T_497 ? tlb_entries_p1_pfn__T_7_data : tlb_entries_p0_pfn__T_7_data; // @[tlb.scala 56:19]
  wire  _T_498_v = _T_497 ? tlb_entries_p1_v__T_7_data : tlb_entries_p0_v__T_7_data; // @[tlb.scala 56:19]
  wire  _T_503 = ~_T_498_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1303 = {{8'd0}, _T_498_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_508 = _GEN_1303 & _T_59; // @[tlb.scala 68:32]
  wire [43:0] _T_509 = {_T_508, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_514 = _T_495 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_515 = _GEN_1296 & _T_514; // @[tlb.scala 69:27]
  wire [43:0] _T_516 = _T_509 | _T_515; // @[tlb.scala 70:29]
  wire [4:0] _GEN_19 = _T_503 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_21 = _T_503 ? 44'h0 : _T_516; // @[tlb.scala 59:27]
  wire [31:0] _T_520 = _T_68 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_521 = {_T_520, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_522 = _GEN_1296 & _T_521; // @[tlb.scala 55:24]
  wire  _T_523 = _T_522 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_524_pfn = _T_523 ? tlb_entries_p1_pfn__T_8_data : tlb_entries_p0_pfn__T_8_data; // @[tlb.scala 56:19]
  wire  _T_524_v = _T_523 ? tlb_entries_p1_v__T_8_data : tlb_entries_p0_v__T_8_data; // @[tlb.scala 56:19]
  wire  _T_529 = ~_T_524_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1306 = {{8'd0}, _T_524_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_534 = _GEN_1306 & _T_69; // @[tlb.scala 68:32]
  wire [43:0] _T_535 = {_T_534, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_540 = _T_521 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_541 = _GEN_1296 & _T_540; // @[tlb.scala 69:27]
  wire [43:0] _T_542 = _T_535 | _T_541; // @[tlb.scala 70:29]
  wire [4:0] _GEN_25 = _T_529 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_27 = _T_529 ? 44'h0 : _T_542; // @[tlb.scala 59:27]
  wire [31:0] _T_546 = _T_78 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_547 = {_T_546, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_548 = _GEN_1296 & _T_547; // @[tlb.scala 55:24]
  wire  _T_549 = _T_548 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_550_pfn = _T_549 ? tlb_entries_p1_pfn__T_9_data : tlb_entries_p0_pfn__T_9_data; // @[tlb.scala 56:19]
  wire  _T_550_v = _T_549 ? tlb_entries_p1_v__T_9_data : tlb_entries_p0_v__T_9_data; // @[tlb.scala 56:19]
  wire  _T_555 = ~_T_550_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1309 = {{8'd0}, _T_550_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_560 = _GEN_1309 & _T_79; // @[tlb.scala 68:32]
  wire [43:0] _T_561 = {_T_560, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_566 = _T_547 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_567 = _GEN_1296 & _T_566; // @[tlb.scala 69:27]
  wire [43:0] _T_568 = _T_561 | _T_567; // @[tlb.scala 70:29]
  wire [4:0] _GEN_31 = _T_555 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_33 = _T_555 ? 44'h0 : _T_568; // @[tlb.scala 59:27]
  wire [31:0] _T_572 = _T_88 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_573 = {_T_572, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_574 = _GEN_1296 & _T_573; // @[tlb.scala 55:24]
  wire  _T_575 = _T_574 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_576_pfn = _T_575 ? tlb_entries_p1_pfn__T_10_data : tlb_entries_p0_pfn__T_10_data; // @[tlb.scala 56:19]
  wire  _T_576_v = _T_575 ? tlb_entries_p1_v__T_10_data : tlb_entries_p0_v__T_10_data; // @[tlb.scala 56:19]
  wire  _T_581 = ~_T_576_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1312 = {{8'd0}, _T_576_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_586 = _GEN_1312 & _T_89; // @[tlb.scala 68:32]
  wire [43:0] _T_587 = {_T_586, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_592 = _T_573 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_593 = _GEN_1296 & _T_592; // @[tlb.scala 69:27]
  wire [43:0] _T_594 = _T_587 | _T_593; // @[tlb.scala 70:29]
  wire [4:0] _GEN_37 = _T_581 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_39 = _T_581 ? 44'h0 : _T_594; // @[tlb.scala 59:27]
  wire [31:0] _T_598 = _T_98 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_599 = {_T_598, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_600 = _GEN_1296 & _T_599; // @[tlb.scala 55:24]
  wire  _T_601 = _T_600 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_602_pfn = _T_601 ? tlb_entries_p1_pfn__T_11_data : tlb_entries_p0_pfn__T_11_data; // @[tlb.scala 56:19]
  wire  _T_602_v = _T_601 ? tlb_entries_p1_v__T_11_data : tlb_entries_p0_v__T_11_data; // @[tlb.scala 56:19]
  wire  _T_607 = ~_T_602_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1315 = {{8'd0}, _T_602_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_612 = _GEN_1315 & _T_99; // @[tlb.scala 68:32]
  wire [43:0] _T_613 = {_T_612, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_618 = _T_599 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_619 = _GEN_1296 & _T_618; // @[tlb.scala 69:27]
  wire [43:0] _T_620 = _T_613 | _T_619; // @[tlb.scala 70:29]
  wire [4:0] _GEN_43 = _T_607 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_45 = _T_607 ? 44'h0 : _T_620; // @[tlb.scala 59:27]
  wire [31:0] _T_624 = _T_108 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_625 = {_T_624, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_626 = _GEN_1296 & _T_625; // @[tlb.scala 55:24]
  wire  _T_627 = _T_626 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_628_pfn = _T_627 ? tlb_entries_p1_pfn__T_12_data : tlb_entries_p0_pfn__T_12_data; // @[tlb.scala 56:19]
  wire  _T_628_v = _T_627 ? tlb_entries_p1_v__T_12_data : tlb_entries_p0_v__T_12_data; // @[tlb.scala 56:19]
  wire  _T_633 = ~_T_628_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1318 = {{8'd0}, _T_628_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_638 = _GEN_1318 & _T_109; // @[tlb.scala 68:32]
  wire [43:0] _T_639 = {_T_638, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_644 = _T_625 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_645 = _GEN_1296 & _T_644; // @[tlb.scala 69:27]
  wire [43:0] _T_646 = _T_639 | _T_645; // @[tlb.scala 70:29]
  wire [4:0] _GEN_49 = _T_633 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_51 = _T_633 ? 44'h0 : _T_646; // @[tlb.scala 59:27]
  wire [31:0] _T_650 = _T_118 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_651 = {_T_650, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_652 = _GEN_1296 & _T_651; // @[tlb.scala 55:24]
  wire  _T_653 = _T_652 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_654_pfn = _T_653 ? tlb_entries_p1_pfn__T_13_data : tlb_entries_p0_pfn__T_13_data; // @[tlb.scala 56:19]
  wire  _T_654_v = _T_653 ? tlb_entries_p1_v__T_13_data : tlb_entries_p0_v__T_13_data; // @[tlb.scala 56:19]
  wire  _T_659 = ~_T_654_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1321 = {{8'd0}, _T_654_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_664 = _GEN_1321 & _T_119; // @[tlb.scala 68:32]
  wire [43:0] _T_665 = {_T_664, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_670 = _T_651 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_671 = _GEN_1296 & _T_670; // @[tlb.scala 69:27]
  wire [43:0] _T_672 = _T_665 | _T_671; // @[tlb.scala 70:29]
  wire [4:0] _GEN_55 = _T_659 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_57 = _T_659 ? 44'h0 : _T_672; // @[tlb.scala 59:27]
  wire [31:0] _T_676 = _T_128 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_677 = {_T_676, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_678 = _GEN_1296 & _T_677; // @[tlb.scala 55:24]
  wire  _T_679 = _T_678 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_680_pfn = _T_679 ? tlb_entries_p1_pfn__T_14_data : tlb_entries_p0_pfn__T_14_data; // @[tlb.scala 56:19]
  wire  _T_680_v = _T_679 ? tlb_entries_p1_v__T_14_data : tlb_entries_p0_v__T_14_data; // @[tlb.scala 56:19]
  wire  _T_685 = ~_T_680_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1324 = {{8'd0}, _T_680_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_690 = _GEN_1324 & _T_129; // @[tlb.scala 68:32]
  wire [43:0] _T_691 = {_T_690, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_696 = _T_677 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_697 = _GEN_1296 & _T_696; // @[tlb.scala 69:27]
  wire [43:0] _T_698 = _T_691 | _T_697; // @[tlb.scala 70:29]
  wire [4:0] _GEN_61 = _T_685 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_63 = _T_685 ? 44'h0 : _T_698; // @[tlb.scala 59:27]
  wire [31:0] _T_702 = _T_138 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_703 = {_T_702, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_704 = _GEN_1296 & _T_703; // @[tlb.scala 55:24]
  wire  _T_705 = _T_704 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_706_pfn = _T_705 ? tlb_entries_p1_pfn__T_15_data : tlb_entries_p0_pfn__T_15_data; // @[tlb.scala 56:19]
  wire  _T_706_v = _T_705 ? tlb_entries_p1_v__T_15_data : tlb_entries_p0_v__T_15_data; // @[tlb.scala 56:19]
  wire  _T_711 = ~_T_706_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1327 = {{8'd0}, _T_706_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_716 = _GEN_1327 & _T_139; // @[tlb.scala 68:32]
  wire [43:0] _T_717 = {_T_716, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_722 = _T_703 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_723 = _GEN_1296 & _T_722; // @[tlb.scala 69:27]
  wire [43:0] _T_724 = _T_717 | _T_723; // @[tlb.scala 70:29]
  wire [4:0] _GEN_67 = _T_711 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_69 = _T_711 ? 44'h0 : _T_724; // @[tlb.scala 59:27]
  wire [31:0] _T_728 = _T_148 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_729 = {_T_728, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_730 = _GEN_1296 & _T_729; // @[tlb.scala 55:24]
  wire  _T_731 = _T_730 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_732_pfn = _T_731 ? tlb_entries_p1_pfn__T_16_data : tlb_entries_p0_pfn__T_16_data; // @[tlb.scala 56:19]
  wire  _T_732_v = _T_731 ? tlb_entries_p1_v__T_16_data : tlb_entries_p0_v__T_16_data; // @[tlb.scala 56:19]
  wire  _T_737 = ~_T_732_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1330 = {{8'd0}, _T_732_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_742 = _GEN_1330 & _T_149; // @[tlb.scala 68:32]
  wire [43:0] _T_743 = {_T_742, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_748 = _T_729 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_749 = _GEN_1296 & _T_748; // @[tlb.scala 69:27]
  wire [43:0] _T_750 = _T_743 | _T_749; // @[tlb.scala 70:29]
  wire [4:0] _GEN_73 = _T_737 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_75 = _T_737 ? 44'h0 : _T_750; // @[tlb.scala 59:27]
  wire [31:0] _T_754 = _T_158 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_755 = {_T_754, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_756 = _GEN_1296 & _T_755; // @[tlb.scala 55:24]
  wire  _T_757 = _T_756 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_758_pfn = _T_757 ? tlb_entries_p1_pfn__T_17_data : tlb_entries_p0_pfn__T_17_data; // @[tlb.scala 56:19]
  wire  _T_758_v = _T_757 ? tlb_entries_p1_v__T_17_data : tlb_entries_p0_v__T_17_data; // @[tlb.scala 56:19]
  wire  _T_763 = ~_T_758_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1333 = {{8'd0}, _T_758_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_768 = _GEN_1333 & _T_159; // @[tlb.scala 68:32]
  wire [43:0] _T_769 = {_T_768, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_774 = _T_755 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_775 = _GEN_1296 & _T_774; // @[tlb.scala 69:27]
  wire [43:0] _T_776 = _T_769 | _T_775; // @[tlb.scala 70:29]
  wire [4:0] _GEN_79 = _T_763 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_81 = _T_763 ? 44'h0 : _T_776; // @[tlb.scala 59:27]
  wire [31:0] _T_780 = _T_168 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_781 = {_T_780, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_782 = _GEN_1296 & _T_781; // @[tlb.scala 55:24]
  wire  _T_783 = _T_782 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_784_pfn = _T_783 ? tlb_entries_p1_pfn__T_18_data : tlb_entries_p0_pfn__T_18_data; // @[tlb.scala 56:19]
  wire  _T_784_v = _T_783 ? tlb_entries_p1_v__T_18_data : tlb_entries_p0_v__T_18_data; // @[tlb.scala 56:19]
  wire  _T_789 = ~_T_784_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1336 = {{8'd0}, _T_784_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_794 = _GEN_1336 & _T_169; // @[tlb.scala 68:32]
  wire [43:0] _T_795 = {_T_794, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_800 = _T_781 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_801 = _GEN_1296 & _T_800; // @[tlb.scala 69:27]
  wire [43:0] _T_802 = _T_795 | _T_801; // @[tlb.scala 70:29]
  wire [4:0] _GEN_85 = _T_789 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_87 = _T_789 ? 44'h0 : _T_802; // @[tlb.scala 59:27]
  wire [31:0] _T_806 = _T_178 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_807 = {_T_806, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_808 = _GEN_1296 & _T_807; // @[tlb.scala 55:24]
  wire  _T_809 = _T_808 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_810_pfn = _T_809 ? tlb_entries_p1_pfn__T_19_data : tlb_entries_p0_pfn__T_19_data; // @[tlb.scala 56:19]
  wire  _T_810_v = _T_809 ? tlb_entries_p1_v__T_19_data : tlb_entries_p0_v__T_19_data; // @[tlb.scala 56:19]
  wire  _T_815 = ~_T_810_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1339 = {{8'd0}, _T_810_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_820 = _GEN_1339 & _T_179; // @[tlb.scala 68:32]
  wire [43:0] _T_821 = {_T_820, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_826 = _T_807 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_827 = _GEN_1296 & _T_826; // @[tlb.scala 69:27]
  wire [43:0] _T_828 = _T_821 | _T_827; // @[tlb.scala 70:29]
  wire [4:0] _GEN_91 = _T_815 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_93 = _T_815 ? 44'h0 : _T_828; // @[tlb.scala 59:27]
  wire [31:0] _T_832 = _T_188 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_833 = {_T_832, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_834 = _GEN_1296 & _T_833; // @[tlb.scala 55:24]
  wire  _T_835 = _T_834 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_836_pfn = _T_835 ? tlb_entries_p1_pfn__T_20_data : tlb_entries_p0_pfn__T_20_data; // @[tlb.scala 56:19]
  wire  _T_836_v = _T_835 ? tlb_entries_p1_v__T_20_data : tlb_entries_p0_v__T_20_data; // @[tlb.scala 56:19]
  wire  _T_841 = ~_T_836_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1342 = {{8'd0}, _T_836_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_846 = _GEN_1342 & _T_189; // @[tlb.scala 68:32]
  wire [43:0] _T_847 = {_T_846, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_852 = _T_833 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_853 = _GEN_1296 & _T_852; // @[tlb.scala 69:27]
  wire [43:0] _T_854 = _T_847 | _T_853; // @[tlb.scala 70:29]
  wire [4:0] _GEN_97 = _T_841 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_99 = _T_841 ? 44'h0 : _T_854; // @[tlb.scala 59:27]
  wire [31:0] _T_858 = _T_198 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_859 = {_T_858, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_860 = _GEN_1296 & _T_859; // @[tlb.scala 55:24]
  wire  _T_861 = _T_860 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_862_pfn = _T_861 ? tlb_entries_p1_pfn__T_21_data : tlb_entries_p0_pfn__T_21_data; // @[tlb.scala 56:19]
  wire  _T_862_v = _T_861 ? tlb_entries_p1_v__T_21_data : tlb_entries_p0_v__T_21_data; // @[tlb.scala 56:19]
  wire  _T_867 = ~_T_862_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1345 = {{8'd0}, _T_862_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_872 = _GEN_1345 & _T_199; // @[tlb.scala 68:32]
  wire [43:0] _T_873 = {_T_872, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_878 = _T_859 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_879 = _GEN_1296 & _T_878; // @[tlb.scala 69:27]
  wire [43:0] _T_880 = _T_873 | _T_879; // @[tlb.scala 70:29]
  wire [4:0] _GEN_103 = _T_867 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_105 = _T_867 ? 44'h0 : _T_880; // @[tlb.scala 59:27]
  wire [31:0] _T_884 = _T_208 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_885 = {_T_884, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_886 = _GEN_1296 & _T_885; // @[tlb.scala 55:24]
  wire  _T_887 = _T_886 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_888_pfn = _T_887 ? tlb_entries_p1_pfn__T_22_data : tlb_entries_p0_pfn__T_22_data; // @[tlb.scala 56:19]
  wire  _T_888_v = _T_887 ? tlb_entries_p1_v__T_22_data : tlb_entries_p0_v__T_22_data; // @[tlb.scala 56:19]
  wire  _T_893 = ~_T_888_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1348 = {{8'd0}, _T_888_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_898 = _GEN_1348 & _T_209; // @[tlb.scala 68:32]
  wire [43:0] _T_899 = {_T_898, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_904 = _T_885 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_905 = _GEN_1296 & _T_904; // @[tlb.scala 69:27]
  wire [43:0] _T_906 = _T_899 | _T_905; // @[tlb.scala 70:29]
  wire [4:0] _GEN_109 = _T_893 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_111 = _T_893 ? 44'h0 : _T_906; // @[tlb.scala 59:27]
  wire [31:0] _T_910 = _T_218 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_911 = {_T_910, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_912 = _GEN_1296 & _T_911; // @[tlb.scala 55:24]
  wire  _T_913 = _T_912 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_914_pfn = _T_913 ? tlb_entries_p1_pfn__T_23_data : tlb_entries_p0_pfn__T_23_data; // @[tlb.scala 56:19]
  wire  _T_914_v = _T_913 ? tlb_entries_p1_v__T_23_data : tlb_entries_p0_v__T_23_data; // @[tlb.scala 56:19]
  wire  _T_919 = ~_T_914_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1351 = {{8'd0}, _T_914_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_924 = _GEN_1351 & _T_219; // @[tlb.scala 68:32]
  wire [43:0] _T_925 = {_T_924, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_930 = _T_911 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_931 = _GEN_1296 & _T_930; // @[tlb.scala 69:27]
  wire [43:0] _T_932 = _T_925 | _T_931; // @[tlb.scala 70:29]
  wire [4:0] _GEN_115 = _T_919 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_117 = _T_919 ? 44'h0 : _T_932; // @[tlb.scala 59:27]
  wire [31:0] _T_936 = _T_228 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_937 = {_T_936, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_938 = _GEN_1296 & _T_937; // @[tlb.scala 55:24]
  wire  _T_939 = _T_938 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_940_pfn = _T_939 ? tlb_entries_p1_pfn__T_24_data : tlb_entries_p0_pfn__T_24_data; // @[tlb.scala 56:19]
  wire  _T_940_v = _T_939 ? tlb_entries_p1_v__T_24_data : tlb_entries_p0_v__T_24_data; // @[tlb.scala 56:19]
  wire  _T_945 = ~_T_940_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1354 = {{8'd0}, _T_940_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_950 = _GEN_1354 & _T_229; // @[tlb.scala 68:32]
  wire [43:0] _T_951 = {_T_950, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_956 = _T_937 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_957 = _GEN_1296 & _T_956; // @[tlb.scala 69:27]
  wire [43:0] _T_958 = _T_951 | _T_957; // @[tlb.scala 70:29]
  wire [4:0] _GEN_121 = _T_945 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_123 = _T_945 ? 44'h0 : _T_958; // @[tlb.scala 59:27]
  wire [31:0] _T_962 = _T_238 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_963 = {_T_962, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_964 = _GEN_1296 & _T_963; // @[tlb.scala 55:24]
  wire  _T_965 = _T_964 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_966_pfn = _T_965 ? tlb_entries_p1_pfn__T_25_data : tlb_entries_p0_pfn__T_25_data; // @[tlb.scala 56:19]
  wire  _T_966_v = _T_965 ? tlb_entries_p1_v__T_25_data : tlb_entries_p0_v__T_25_data; // @[tlb.scala 56:19]
  wire  _T_971 = ~_T_966_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1357 = {{8'd0}, _T_966_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_976 = _GEN_1357 & _T_239; // @[tlb.scala 68:32]
  wire [43:0] _T_977 = {_T_976, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_982 = _T_963 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_983 = _GEN_1296 & _T_982; // @[tlb.scala 69:27]
  wire [43:0] _T_984 = _T_977 | _T_983; // @[tlb.scala 70:29]
  wire [4:0] _GEN_127 = _T_971 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_129 = _T_971 ? 44'h0 : _T_984; // @[tlb.scala 59:27]
  wire [31:0] _T_988 = _T_248 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_989 = {_T_988, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_990 = _GEN_1296 & _T_989; // @[tlb.scala 55:24]
  wire  _T_991 = _T_990 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_992_pfn = _T_991 ? tlb_entries_p1_pfn__T_26_data : tlb_entries_p0_pfn__T_26_data; // @[tlb.scala 56:19]
  wire  _T_992_v = _T_991 ? tlb_entries_p1_v__T_26_data : tlb_entries_p0_v__T_26_data; // @[tlb.scala 56:19]
  wire  _T_997 = ~_T_992_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1360 = {{8'd0}, _T_992_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1002 = _GEN_1360 & _T_249; // @[tlb.scala 68:32]
  wire [43:0] _T_1003 = {_T_1002, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1008 = _T_989 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1009 = _GEN_1296 & _T_1008; // @[tlb.scala 69:27]
  wire [43:0] _T_1010 = _T_1003 | _T_1009; // @[tlb.scala 70:29]
  wire [4:0] _GEN_133 = _T_997 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_135 = _T_997 ? 44'h0 : _T_1010; // @[tlb.scala 59:27]
  wire [31:0] _T_1014 = _T_258 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1015 = {_T_1014, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1016 = _GEN_1296 & _T_1015; // @[tlb.scala 55:24]
  wire  _T_1017 = _T_1016 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1018_pfn = _T_1017 ? tlb_entries_p1_pfn__T_27_data : tlb_entries_p0_pfn__T_27_data; // @[tlb.scala 56:19]
  wire  _T_1018_v = _T_1017 ? tlb_entries_p1_v__T_27_data : tlb_entries_p0_v__T_27_data; // @[tlb.scala 56:19]
  wire  _T_1023 = ~_T_1018_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1363 = {{8'd0}, _T_1018_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1028 = _GEN_1363 & _T_259; // @[tlb.scala 68:32]
  wire [43:0] _T_1029 = {_T_1028, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1034 = _T_1015 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1035 = _GEN_1296 & _T_1034; // @[tlb.scala 69:27]
  wire [43:0] _T_1036 = _T_1029 | _T_1035; // @[tlb.scala 70:29]
  wire [4:0] _GEN_139 = _T_1023 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_141 = _T_1023 ? 44'h0 : _T_1036; // @[tlb.scala 59:27]
  wire [31:0] _T_1040 = _T_268 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1041 = {_T_1040, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1042 = _GEN_1296 & _T_1041; // @[tlb.scala 55:24]
  wire  _T_1043 = _T_1042 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1044_pfn = _T_1043 ? tlb_entries_p1_pfn__T_28_data : tlb_entries_p0_pfn__T_28_data; // @[tlb.scala 56:19]
  wire  _T_1044_v = _T_1043 ? tlb_entries_p1_v__T_28_data : tlb_entries_p0_v__T_28_data; // @[tlb.scala 56:19]
  wire  _T_1049 = ~_T_1044_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1366 = {{8'd0}, _T_1044_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1054 = _GEN_1366 & _T_269; // @[tlb.scala 68:32]
  wire [43:0] _T_1055 = {_T_1054, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1060 = _T_1041 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1061 = _GEN_1296 & _T_1060; // @[tlb.scala 69:27]
  wire [43:0] _T_1062 = _T_1055 | _T_1061; // @[tlb.scala 70:29]
  wire [4:0] _GEN_145 = _T_1049 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_147 = _T_1049 ? 44'h0 : _T_1062; // @[tlb.scala 59:27]
  wire [31:0] _T_1066 = _T_278 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1067 = {_T_1066, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1068 = _GEN_1296 & _T_1067; // @[tlb.scala 55:24]
  wire  _T_1069 = _T_1068 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1070_pfn = _T_1069 ? tlb_entries_p1_pfn__T_29_data : tlb_entries_p0_pfn__T_29_data; // @[tlb.scala 56:19]
  wire  _T_1070_v = _T_1069 ? tlb_entries_p1_v__T_29_data : tlb_entries_p0_v__T_29_data; // @[tlb.scala 56:19]
  wire  _T_1075 = ~_T_1070_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1369 = {{8'd0}, _T_1070_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1080 = _GEN_1369 & _T_279; // @[tlb.scala 68:32]
  wire [43:0] _T_1081 = {_T_1080, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1086 = _T_1067 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1087 = _GEN_1296 & _T_1086; // @[tlb.scala 69:27]
  wire [43:0] _T_1088 = _T_1081 | _T_1087; // @[tlb.scala 70:29]
  wire [4:0] _GEN_151 = _T_1075 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_153 = _T_1075 ? 44'h0 : _T_1088; // @[tlb.scala 59:27]
  wire [31:0] _T_1092 = _T_288 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1093 = {_T_1092, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1094 = _GEN_1296 & _T_1093; // @[tlb.scala 55:24]
  wire  _T_1095 = _T_1094 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1096_pfn = _T_1095 ? tlb_entries_p1_pfn__T_30_data : tlb_entries_p0_pfn__T_30_data; // @[tlb.scala 56:19]
  wire  _T_1096_v = _T_1095 ? tlb_entries_p1_v__T_30_data : tlb_entries_p0_v__T_30_data; // @[tlb.scala 56:19]
  wire  _T_1101 = ~_T_1096_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1372 = {{8'd0}, _T_1096_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1106 = _GEN_1372 & _T_289; // @[tlb.scala 68:32]
  wire [43:0] _T_1107 = {_T_1106, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1112 = _T_1093 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1113 = _GEN_1296 & _T_1112; // @[tlb.scala 69:27]
  wire [43:0] _T_1114 = _T_1107 | _T_1113; // @[tlb.scala 70:29]
  wire [4:0] _GEN_157 = _T_1101 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_159 = _T_1101 ? 44'h0 : _T_1114; // @[tlb.scala 59:27]
  wire [31:0] _T_1118 = _T_298 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1119 = {_T_1118, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1120 = _GEN_1296 & _T_1119; // @[tlb.scala 55:24]
  wire  _T_1121 = _T_1120 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1122_pfn = _T_1121 ? tlb_entries_p1_pfn__T_31_data : tlb_entries_p0_pfn__T_31_data; // @[tlb.scala 56:19]
  wire  _T_1122_v = _T_1121 ? tlb_entries_p1_v__T_31_data : tlb_entries_p0_v__T_31_data; // @[tlb.scala 56:19]
  wire  _T_1127 = ~_T_1122_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1375 = {{8'd0}, _T_1122_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1132 = _GEN_1375 & _T_299; // @[tlb.scala 68:32]
  wire [43:0] _T_1133 = {_T_1132, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1138 = _T_1119 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1139 = _GEN_1296 & _T_1138; // @[tlb.scala 69:27]
  wire [43:0] _T_1140 = _T_1133 | _T_1139; // @[tlb.scala 70:29]
  wire [4:0] _GEN_163 = _T_1127 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_165 = _T_1127 ? 44'h0 : _T_1140; // @[tlb.scala 59:27]
  wire [31:0] _T_1144 = _T_308 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1145 = {_T_1144, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1146 = _GEN_1296 & _T_1145; // @[tlb.scala 55:24]
  wire  _T_1147 = _T_1146 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1148_pfn = _T_1147 ? tlb_entries_p1_pfn__T_32_data : tlb_entries_p0_pfn__T_32_data; // @[tlb.scala 56:19]
  wire  _T_1148_v = _T_1147 ? tlb_entries_p1_v__T_32_data : tlb_entries_p0_v__T_32_data; // @[tlb.scala 56:19]
  wire  _T_1153 = ~_T_1148_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1378 = {{8'd0}, _T_1148_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1158 = _GEN_1378 & _T_309; // @[tlb.scala 68:32]
  wire [43:0] _T_1159 = {_T_1158, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1164 = _T_1145 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1165 = _GEN_1296 & _T_1164; // @[tlb.scala 69:27]
  wire [43:0] _T_1166 = _T_1159 | _T_1165; // @[tlb.scala 70:29]
  wire [4:0] _GEN_169 = _T_1153 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_171 = _T_1153 ? 44'h0 : _T_1166; // @[tlb.scala 59:27]
  wire [31:0] _T_1170 = _T_318 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1171 = {_T_1170, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1172 = _GEN_1296 & _T_1171; // @[tlb.scala 55:24]
  wire  _T_1173 = _T_1172 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1174_pfn = _T_1173 ? tlb_entries_p1_pfn__T_33_data : tlb_entries_p0_pfn__T_33_data; // @[tlb.scala 56:19]
  wire  _T_1174_v = _T_1173 ? tlb_entries_p1_v__T_33_data : tlb_entries_p0_v__T_33_data; // @[tlb.scala 56:19]
  wire  _T_1179 = ~_T_1174_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1381 = {{8'd0}, _T_1174_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1184 = _GEN_1381 & _T_319; // @[tlb.scala 68:32]
  wire [43:0] _T_1185 = {_T_1184, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1190 = _T_1171 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1191 = _GEN_1296 & _T_1190; // @[tlb.scala 69:27]
  wire [43:0] _T_1192 = _T_1185 | _T_1191; // @[tlb.scala 70:29]
  wire [4:0] _GEN_175 = _T_1179 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_177 = _T_1179 ? 44'h0 : _T_1192; // @[tlb.scala 59:27]
  wire [31:0] _T_1196 = _T_328 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1197 = {_T_1196, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1198 = _GEN_1296 & _T_1197; // @[tlb.scala 55:24]
  wire  _T_1199 = _T_1198 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1200_pfn = _T_1199 ? tlb_entries_p1_pfn__T_34_data : tlb_entries_p0_pfn__T_34_data; // @[tlb.scala 56:19]
  wire  _T_1200_v = _T_1199 ? tlb_entries_p1_v__T_34_data : tlb_entries_p0_v__T_34_data; // @[tlb.scala 56:19]
  wire  _T_1205 = ~_T_1200_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1384 = {{8'd0}, _T_1200_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1210 = _GEN_1384 & _T_329; // @[tlb.scala 68:32]
  wire [43:0] _T_1211 = {_T_1210, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1216 = _T_1197 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1217 = _GEN_1296 & _T_1216; // @[tlb.scala 69:27]
  wire [43:0] _T_1218 = _T_1211 | _T_1217; // @[tlb.scala 70:29]
  wire [4:0] _GEN_181 = _T_1205 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_183 = _T_1205 ? 44'h0 : _T_1218; // @[tlb.scala 59:27]
  wire [31:0] _T_1222 = _T_338 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1223 = {_T_1222, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1224 = _GEN_1296 & _T_1223; // @[tlb.scala 55:24]
  wire  _T_1225 = _T_1224 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1226_pfn = _T_1225 ? tlb_entries_p1_pfn__T_35_data : tlb_entries_p0_pfn__T_35_data; // @[tlb.scala 56:19]
  wire  _T_1226_v = _T_1225 ? tlb_entries_p1_v__T_35_data : tlb_entries_p0_v__T_35_data; // @[tlb.scala 56:19]
  wire  _T_1231 = ~_T_1226_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1387 = {{8'd0}, _T_1226_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1236 = _GEN_1387 & _T_339; // @[tlb.scala 68:32]
  wire [43:0] _T_1237 = {_T_1236, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1242 = _T_1223 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1243 = _GEN_1296 & _T_1242; // @[tlb.scala 69:27]
  wire [43:0] _T_1244 = _T_1237 | _T_1243; // @[tlb.scala 70:29]
  wire [4:0] _GEN_187 = _T_1231 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_189 = _T_1231 ? 44'h0 : _T_1244; // @[tlb.scala 59:27]
  wire [31:0] _T_1248 = _T_348 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1249 = {_T_1248, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_1250 = _GEN_1296 & _T_1249; // @[tlb.scala 55:24]
  wire  _T_1251 = _T_1250 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1252_pfn = _T_1251 ? tlb_entries_p1_pfn__T_36_data : tlb_entries_p0_pfn__T_36_data; // @[tlb.scala 56:19]
  wire  _T_1252_v = _T_1251 ? tlb_entries_p1_v__T_36_data : tlb_entries_p0_v__T_36_data; // @[tlb.scala 56:19]
  wire  _T_1257 = ~_T_1252_v; // @[tlb.scala 59:18]
  wire [31:0] _GEN_1390 = {{8'd0}, _T_1252_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1262 = _GEN_1390 & _T_349; // @[tlb.scala 68:32]
  wire [43:0] _T_1263 = {_T_1262, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_1268 = _T_1249 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_1269 = _GEN_1296 & _T_1268; // @[tlb.scala 69:27]
  wire [43:0] _T_1270 = _T_1263 | _T_1269; // @[tlb.scala 70:29]
  wire [4:0] _GEN_193 = _T_1257 ? 5'h8 : 5'h0; // @[tlb.scala 59:27]
  wire [43:0] _GEN_195 = _T_1257 ? 44'h0 : _T_1270; // @[tlb.scala 59:27]
  wire [7:0] _T_450_ex_asid = tlb_entries_asid__T_5_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1274 = {_GEN_7,5'h2,_T_3_vaddr,_T_450_ex_asid,_GEN_9[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1275 = _T_436[0] ? _T_1274 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_476_ex_asid = tlb_entries_asid__T_6_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1279 = {_GEN_13,5'h2,_T_3_vaddr,_T_476_ex_asid,_GEN_15[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1280 = _T_436[1] ? _T_1279 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_502_ex_asid = tlb_entries_asid__T_7_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1284 = {_GEN_19,5'h2,_T_3_vaddr,_T_502_ex_asid,_GEN_21[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1285 = _T_436[2] ? _T_1284 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_528_ex_asid = tlb_entries_asid__T_8_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1289 = {_GEN_25,5'h2,_T_3_vaddr,_T_528_ex_asid,_GEN_27[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1290 = _T_436[3] ? _T_1289 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_554_ex_asid = tlb_entries_asid__T_9_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1294 = {_GEN_31,5'h2,_T_3_vaddr,_T_554_ex_asid,_GEN_33[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1295 = _T_436[4] ? _T_1294 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_580_ex_asid = tlb_entries_asid__T_10_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1299 = {_GEN_37,5'h2,_T_3_vaddr,_T_580_ex_asid,_GEN_39[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1300 = _T_436[5] ? _T_1299 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_606_ex_asid = tlb_entries_asid__T_11_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1304 = {_GEN_43,5'h2,_T_3_vaddr,_T_606_ex_asid,_GEN_45[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1305 = _T_436[6] ? _T_1304 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_632_ex_asid = tlb_entries_asid__T_12_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1309 = {_GEN_49,5'h2,_T_3_vaddr,_T_632_ex_asid,_GEN_51[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1310 = _T_436[7] ? _T_1309 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_658_ex_asid = tlb_entries_asid__T_13_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1314 = {_GEN_55,5'h2,_T_3_vaddr,_T_658_ex_asid,_GEN_57[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1315 = _T_436[8] ? _T_1314 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_684_ex_asid = tlb_entries_asid__T_14_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1319 = {_GEN_61,5'h2,_T_3_vaddr,_T_684_ex_asid,_GEN_63[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1320 = _T_436[9] ? _T_1319 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_710_ex_asid = tlb_entries_asid__T_15_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1324 = {_GEN_67,5'h2,_T_3_vaddr,_T_710_ex_asid,_GEN_69[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1325 = _T_436[10] ? _T_1324 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_736_ex_asid = tlb_entries_asid__T_16_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1329 = {_GEN_73,5'h2,_T_3_vaddr,_T_736_ex_asid,_GEN_75[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1330 = _T_436[11] ? _T_1329 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_762_ex_asid = tlb_entries_asid__T_17_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1334 = {_GEN_79,5'h2,_T_3_vaddr,_T_762_ex_asid,_GEN_81[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1335 = _T_436[12] ? _T_1334 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_788_ex_asid = tlb_entries_asid__T_18_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1339 = {_GEN_85,5'h2,_T_3_vaddr,_T_788_ex_asid,_GEN_87[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1340 = _T_436[13] ? _T_1339 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_814_ex_asid = tlb_entries_asid__T_19_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1344 = {_GEN_91,5'h2,_T_3_vaddr,_T_814_ex_asid,_GEN_93[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1345 = _T_436[14] ? _T_1344 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_840_ex_asid = tlb_entries_asid__T_20_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1349 = {_GEN_97,5'h2,_T_3_vaddr,_T_840_ex_asid,_GEN_99[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1350 = _T_436[15] ? _T_1349 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_866_ex_asid = tlb_entries_asid__T_21_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1354 = {_GEN_103,5'h2,_T_3_vaddr,_T_866_ex_asid,_GEN_105[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1355 = _T_436[16] ? _T_1354 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_892_ex_asid = tlb_entries_asid__T_22_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1359 = {_GEN_109,5'h2,_T_3_vaddr,_T_892_ex_asid,_GEN_111[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1360 = _T_436[17] ? _T_1359 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_918_ex_asid = tlb_entries_asid__T_23_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1364 = {_GEN_115,5'h2,_T_3_vaddr,_T_918_ex_asid,_GEN_117[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1365 = _T_436[18] ? _T_1364 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_944_ex_asid = tlb_entries_asid__T_24_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1369 = {_GEN_121,5'h2,_T_3_vaddr,_T_944_ex_asid,_GEN_123[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1370 = _T_436[19] ? _T_1369 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_970_ex_asid = tlb_entries_asid__T_25_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1374 = {_GEN_127,5'h2,_T_3_vaddr,_T_970_ex_asid,_GEN_129[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1375 = _T_436[20] ? _T_1374 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_996_ex_asid = tlb_entries_asid__T_26_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1379 = {_GEN_133,5'h2,_T_3_vaddr,_T_996_ex_asid,_GEN_135[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1380 = _T_436[21] ? _T_1379 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1022_ex_asid = tlb_entries_asid__T_27_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1384 = {_GEN_139,5'h2,_T_3_vaddr,_T_1022_ex_asid,_GEN_141[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1385 = _T_436[22] ? _T_1384 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1048_ex_asid = tlb_entries_asid__T_28_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1389 = {_GEN_145,5'h2,_T_3_vaddr,_T_1048_ex_asid,_GEN_147[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1390 = _T_436[23] ? _T_1389 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1074_ex_asid = tlb_entries_asid__T_29_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1394 = {_GEN_151,5'h2,_T_3_vaddr,_T_1074_ex_asid,_GEN_153[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1395 = _T_436[24] ? _T_1394 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1100_ex_asid = tlb_entries_asid__T_30_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1399 = {_GEN_157,5'h2,_T_3_vaddr,_T_1100_ex_asid,_GEN_159[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1400 = _T_436[25] ? _T_1399 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1126_ex_asid = tlb_entries_asid__T_31_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1404 = {_GEN_163,5'h2,_T_3_vaddr,_T_1126_ex_asid,_GEN_165[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1405 = _T_436[26] ? _T_1404 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1152_ex_asid = tlb_entries_asid__T_32_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1409 = {_GEN_169,5'h2,_T_3_vaddr,_T_1152_ex_asid,_GEN_171[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1410 = _T_436[27] ? _T_1409 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1178_ex_asid = tlb_entries_asid__T_33_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1414 = {_GEN_175,5'h2,_T_3_vaddr,_T_1178_ex_asid,_GEN_177[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1415 = _T_436[28] ? _T_1414 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1204_ex_asid = tlb_entries_asid__T_34_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1419 = {_GEN_181,5'h2,_T_3_vaddr,_T_1204_ex_asid,_GEN_183[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1420 = _T_436[29] ? _T_1419 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1230_ex_asid = tlb_entries_asid__T_35_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1424 = {_GEN_187,5'h2,_T_3_vaddr,_T_1230_ex_asid,_GEN_189[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1425 = _T_436[30] ? _T_1424 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1256_ex_asid = tlb_entries_asid__T_36_data; // @[tlb.scala 74:17]
  wire [81:0] _T_1429 = {_GEN_193,5'h2,_T_3_vaddr,_T_1256_ex_asid,_GEN_195[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_1430 = _T_436[31] ? _T_1429 : 82'h0; // @[Mux.scala 27:72]
  wire [81:0] _T_1431 = _T_1275 | _T_1280; // @[Mux.scala 27:72]
  wire [81:0] _T_1432 = _T_1431 | _T_1285; // @[Mux.scala 27:72]
  wire [81:0] _T_1433 = _T_1432 | _T_1290; // @[Mux.scala 27:72]
  wire [81:0] _T_1434 = _T_1433 | _T_1295; // @[Mux.scala 27:72]
  wire [81:0] _T_1435 = _T_1434 | _T_1300; // @[Mux.scala 27:72]
  wire [81:0] _T_1436 = _T_1435 | _T_1305; // @[Mux.scala 27:72]
  wire [81:0] _T_1437 = _T_1436 | _T_1310; // @[Mux.scala 27:72]
  wire [81:0] _T_1438 = _T_1437 | _T_1315; // @[Mux.scala 27:72]
  wire [81:0] _T_1439 = _T_1438 | _T_1320; // @[Mux.scala 27:72]
  wire [81:0] _T_1440 = _T_1439 | _T_1325; // @[Mux.scala 27:72]
  wire [81:0] _T_1441 = _T_1440 | _T_1330; // @[Mux.scala 27:72]
  wire [81:0] _T_1442 = _T_1441 | _T_1335; // @[Mux.scala 27:72]
  wire [81:0] _T_1443 = _T_1442 | _T_1340; // @[Mux.scala 27:72]
  wire [81:0] _T_1444 = _T_1443 | _T_1345; // @[Mux.scala 27:72]
  wire [81:0] _T_1445 = _T_1444 | _T_1350; // @[Mux.scala 27:72]
  wire [81:0] _T_1446 = _T_1445 | _T_1355; // @[Mux.scala 27:72]
  wire [81:0] _T_1447 = _T_1446 | _T_1360; // @[Mux.scala 27:72]
  wire [81:0] _T_1448 = _T_1447 | _T_1365; // @[Mux.scala 27:72]
  wire [81:0] _T_1449 = _T_1448 | _T_1370; // @[Mux.scala 27:72]
  wire [81:0] _T_1450 = _T_1449 | _T_1375; // @[Mux.scala 27:72]
  wire [81:0] _T_1451 = _T_1450 | _T_1380; // @[Mux.scala 27:72]
  wire [81:0] _T_1452 = _T_1451 | _T_1385; // @[Mux.scala 27:72]
  wire [81:0] _T_1453 = _T_1452 | _T_1390; // @[Mux.scala 27:72]
  wire [81:0] _T_1454 = _T_1453 | _T_1395; // @[Mux.scala 27:72]
  wire [81:0] _T_1455 = _T_1454 | _T_1400; // @[Mux.scala 27:72]
  wire [81:0] _T_1456 = _T_1455 | _T_1405; // @[Mux.scala 27:72]
  wire [81:0] _T_1457 = _T_1456 | _T_1410; // @[Mux.scala 27:72]
  wire [81:0] _T_1458 = _T_1457 | _T_1415; // @[Mux.scala 27:72]
  wire [81:0] _T_1459 = _T_1458 | _T_1420; // @[Mux.scala 27:72]
  wire [81:0] _T_1460 = _T_1459 | _T_1425; // @[Mux.scala 27:72]
  wire [81:0] _T_1461 = _T_1460 | _T_1430; // @[Mux.scala 27:72]
  wire [4:0] _T_1473_ex_et = _T_438 ? 5'h7 : _T_1461[81:77]; // @[tlb.scala 102:8]
  wire [4:0] _T_1473_ex_code = _T_438 ? 5'h2 : _T_1461[76:72]; // @[tlb.scala 102:8]
  wire [7:0] _T_1473_ex_asid = _T_438 ? 8'h0 : _T_1461[39:32]; // @[tlb.scala 102:8]
  wire [31:0] _T_1473_paddr = _T_438 ? 32'h0 : _T_1461[31:0]; // @[tlb.scala 102:8]
  wire  _T_1475 = _T_3_vaddr[31:29] == 3'h4; // @[tlb.scala 111:12]
  wire  _T_1476 = _T_3_vaddr[31:29] == 3'h5; // @[tlb.scala 111:27]
  wire  _T_1477 = _T_1475 | _T_1476; // @[tlb.scala 111:20]
  wire [29:0] _T_1479 = {1'h0,_T_3_vaddr[28:0]}; // @[Cat.scala 29:58]
  wire  _T_1480 = _T_3_vaddr[31:29] == 3'h6; // @[tlb.scala 112:12]
  wire [29:0] _T_1482 = {1'h0,_T_1473_paddr[28:0]}; // @[Cat.scala 29:58]
  wire  _T_1483 = _T_3_vaddr[31:29] == 3'h7; // @[tlb.scala 113:12]
  wire  _T_1485 = ~_T_3_vaddr[31]; // @[tlb.scala 114:15]
  wire [31:0] _T_1488 = io_status_ERL ? _T_3_vaddr : {{2'd0}, _T_1482}; // @[tlb.scala 114:30]
  wire [29:0] _T_1489 = _T_1477 ? _T_1479 : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_1490 = _T_1480 ? _T_1482 : 30'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1491 = _T_1483 ? _T_3_vaddr : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1492 = _T_1485 ? _T_1488 : 32'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_1493 = _T_1489 | _T_1490; // @[Mux.scala 27:72]
  wire [31:0] _GEN_1392 = {{2'd0}, _T_1493}; // @[Mux.scala 27:72]
  wire [31:0] _T_1494 = _GEN_1392 | _T_1491; // @[Mux.scala 27:72]
  wire [4:0] _T_1503 = io_status_ERL ? 5'h0 : _T_1473_ex_et; // @[tlb.scala 120:30]
  wire [4:0] _T_1505 = _T_1480 ? _T_1473_ex_et : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1506 = _T_1485 ? _T_1503 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1508 = _T_1505 | _T_1506; // @[Mux.scala 27:72]
  wire [1:0] _T_1513 = _T_3_is_aligned ? _T_3_vaddr[1:0] : 2'h0; // @[tlb.scala 148:23]
  wire  _T_1515 = _T_3_len == 2'h1; // @[tlb.scala 152:22]
  wire  _T_1517 = _T_3_len == 2'h3; // @[tlb.scala 153:22]
  wire  _T_1518 = _T_1513 != 2'h0; // @[tlb.scala 153:45]
  wire  _T_1520 = _T_1515 & _T_1513[0]; // @[Mux.scala 27:72]
  wire  _T_1521 = _T_1517 & _T_1518; // @[Mux.scala 27:72]
  wire  _T_1523 = _T_1520 | _T_1521; // @[Mux.scala 27:72]
  wire  _T_1529 = ~_T_4; // @[tlb.scala 160:40]
  wire  _T_1535 = ~_T_1; // @[tlb.scala 166:21]
  wire  _T_1536 = io_iaddr_resp_ready & io_iaddr_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_1537 = _T_1535 & _T_1536; // @[tlb.scala 166:37]
  wire  _T_1538 = _T | _T_1537; // @[tlb.scala 166:17]
  wire  _T_1539 = ~_T; // @[tlb.scala 168:18]
  wire  _T_1541 = _T_1539 & _T_1; // @[tlb.scala 168:25]
  wire  _GEN_196 = _T_1541 | _T_4; // @[tlb.scala 168:44]
  wire  _T_1542 = io_daddr_req_ready & io_daddr_req_valid; // @[Decoupled.scala 40:37]
  reg  _T_1544_func; // @[Reg.scala 27:20]
  reg [31:0] _RAND_16;
  reg [31:0] _T_1544_vaddr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_17;
  reg [1:0] _T_1544_len; // @[Reg.scala 27:20]
  reg [31:0] _RAND_18;
  reg  _T_1544_is_aligned; // @[Reg.scala 27:20]
  reg [31:0] _RAND_19;
  wire [31:0] _T_1579 = {{16'd0}, tlb_entries_pagemask__T_1546_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1580 = ~_T_1579; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1393 = {{13'd0}, tlb_entries_vpn__T_1546_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1581 = _GEN_1393 & _T_1580; // @[tlb.scala 50:19]
  wire [31:0] _GEN_1394 = {{13'd0}, _T_1544_vaddr[31:13]}; // @[tlb.scala 50:37]
  wire [31:0] _T_1583 = _GEN_1394 & _T_1580; // @[tlb.scala 50:37]
  wire  _T_1584 = _T_1581 == _T_1583; // @[tlb.scala 50:28]
  wire  _T_1585 = tlb_entries_asid__T_1546_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1586 = tlb_entries_g__T_1546_data | _T_1585; // @[tlb.scala 51:17]
  wire  _T_1587 = _T_1584 & _T_1586; // @[tlb.scala 50:46]
  wire [31:0] _T_1589 = {{16'd0}, tlb_entries_pagemask__T_1547_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1590 = ~_T_1589; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1395 = {{13'd0}, tlb_entries_vpn__T_1547_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1591 = _GEN_1395 & _T_1590; // @[tlb.scala 50:19]
  wire [31:0] _T_1593 = _GEN_1394 & _T_1590; // @[tlb.scala 50:37]
  wire  _T_1594 = _T_1591 == _T_1593; // @[tlb.scala 50:28]
  wire  _T_1595 = tlb_entries_asid__T_1547_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1596 = tlb_entries_g__T_1547_data | _T_1595; // @[tlb.scala 51:17]
  wire  _T_1597 = _T_1594 & _T_1596; // @[tlb.scala 50:46]
  wire [31:0] _T_1599 = {{16'd0}, tlb_entries_pagemask__T_1548_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1600 = ~_T_1599; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1397 = {{13'd0}, tlb_entries_vpn__T_1548_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1601 = _GEN_1397 & _T_1600; // @[tlb.scala 50:19]
  wire [31:0] _T_1603 = _GEN_1394 & _T_1600; // @[tlb.scala 50:37]
  wire  _T_1604 = _T_1601 == _T_1603; // @[tlb.scala 50:28]
  wire  _T_1605 = tlb_entries_asid__T_1548_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1606 = tlb_entries_g__T_1548_data | _T_1605; // @[tlb.scala 51:17]
  wire  _T_1607 = _T_1604 & _T_1606; // @[tlb.scala 50:46]
  wire [31:0] _T_1609 = {{16'd0}, tlb_entries_pagemask__T_1549_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1610 = ~_T_1609; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1399 = {{13'd0}, tlb_entries_vpn__T_1549_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1611 = _GEN_1399 & _T_1610; // @[tlb.scala 50:19]
  wire [31:0] _T_1613 = _GEN_1394 & _T_1610; // @[tlb.scala 50:37]
  wire  _T_1614 = _T_1611 == _T_1613; // @[tlb.scala 50:28]
  wire  _T_1615 = tlb_entries_asid__T_1549_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1616 = tlb_entries_g__T_1549_data | _T_1615; // @[tlb.scala 51:17]
  wire  _T_1617 = _T_1614 & _T_1616; // @[tlb.scala 50:46]
  wire [31:0] _T_1619 = {{16'd0}, tlb_entries_pagemask__T_1550_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1620 = ~_T_1619; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1401 = {{13'd0}, tlb_entries_vpn__T_1550_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1621 = _GEN_1401 & _T_1620; // @[tlb.scala 50:19]
  wire [31:0] _T_1623 = _GEN_1394 & _T_1620; // @[tlb.scala 50:37]
  wire  _T_1624 = _T_1621 == _T_1623; // @[tlb.scala 50:28]
  wire  _T_1625 = tlb_entries_asid__T_1550_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1626 = tlb_entries_g__T_1550_data | _T_1625; // @[tlb.scala 51:17]
  wire  _T_1627 = _T_1624 & _T_1626; // @[tlb.scala 50:46]
  wire [31:0] _T_1629 = {{16'd0}, tlb_entries_pagemask__T_1551_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1630 = ~_T_1629; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1403 = {{13'd0}, tlb_entries_vpn__T_1551_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1631 = _GEN_1403 & _T_1630; // @[tlb.scala 50:19]
  wire [31:0] _T_1633 = _GEN_1394 & _T_1630; // @[tlb.scala 50:37]
  wire  _T_1634 = _T_1631 == _T_1633; // @[tlb.scala 50:28]
  wire  _T_1635 = tlb_entries_asid__T_1551_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1636 = tlb_entries_g__T_1551_data | _T_1635; // @[tlb.scala 51:17]
  wire  _T_1637 = _T_1634 & _T_1636; // @[tlb.scala 50:46]
  wire [31:0] _T_1639 = {{16'd0}, tlb_entries_pagemask__T_1552_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1640 = ~_T_1639; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1405 = {{13'd0}, tlb_entries_vpn__T_1552_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1641 = _GEN_1405 & _T_1640; // @[tlb.scala 50:19]
  wire [31:0] _T_1643 = _GEN_1394 & _T_1640; // @[tlb.scala 50:37]
  wire  _T_1644 = _T_1641 == _T_1643; // @[tlb.scala 50:28]
  wire  _T_1645 = tlb_entries_asid__T_1552_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1646 = tlb_entries_g__T_1552_data | _T_1645; // @[tlb.scala 51:17]
  wire  _T_1647 = _T_1644 & _T_1646; // @[tlb.scala 50:46]
  wire [31:0] _T_1649 = {{16'd0}, tlb_entries_pagemask__T_1553_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1650 = ~_T_1649; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1407 = {{13'd0}, tlb_entries_vpn__T_1553_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1651 = _GEN_1407 & _T_1650; // @[tlb.scala 50:19]
  wire [31:0] _T_1653 = _GEN_1394 & _T_1650; // @[tlb.scala 50:37]
  wire  _T_1654 = _T_1651 == _T_1653; // @[tlb.scala 50:28]
  wire  _T_1655 = tlb_entries_asid__T_1553_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1656 = tlb_entries_g__T_1553_data | _T_1655; // @[tlb.scala 51:17]
  wire  _T_1657 = _T_1654 & _T_1656; // @[tlb.scala 50:46]
  wire [31:0] _T_1659 = {{16'd0}, tlb_entries_pagemask__T_1554_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1660 = ~_T_1659; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1409 = {{13'd0}, tlb_entries_vpn__T_1554_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1661 = _GEN_1409 & _T_1660; // @[tlb.scala 50:19]
  wire [31:0] _T_1663 = _GEN_1394 & _T_1660; // @[tlb.scala 50:37]
  wire  _T_1664 = _T_1661 == _T_1663; // @[tlb.scala 50:28]
  wire  _T_1665 = tlb_entries_asid__T_1554_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1666 = tlb_entries_g__T_1554_data | _T_1665; // @[tlb.scala 51:17]
  wire  _T_1667 = _T_1664 & _T_1666; // @[tlb.scala 50:46]
  wire [31:0] _T_1669 = {{16'd0}, tlb_entries_pagemask__T_1555_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1670 = ~_T_1669; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1411 = {{13'd0}, tlb_entries_vpn__T_1555_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1671 = _GEN_1411 & _T_1670; // @[tlb.scala 50:19]
  wire [31:0] _T_1673 = _GEN_1394 & _T_1670; // @[tlb.scala 50:37]
  wire  _T_1674 = _T_1671 == _T_1673; // @[tlb.scala 50:28]
  wire  _T_1675 = tlb_entries_asid__T_1555_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1676 = tlb_entries_g__T_1555_data | _T_1675; // @[tlb.scala 51:17]
  wire  _T_1677 = _T_1674 & _T_1676; // @[tlb.scala 50:46]
  wire [31:0] _T_1679 = {{16'd0}, tlb_entries_pagemask__T_1556_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1680 = ~_T_1679; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1413 = {{13'd0}, tlb_entries_vpn__T_1556_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1681 = _GEN_1413 & _T_1680; // @[tlb.scala 50:19]
  wire [31:0] _T_1683 = _GEN_1394 & _T_1680; // @[tlb.scala 50:37]
  wire  _T_1684 = _T_1681 == _T_1683; // @[tlb.scala 50:28]
  wire  _T_1685 = tlb_entries_asid__T_1556_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1686 = tlb_entries_g__T_1556_data | _T_1685; // @[tlb.scala 51:17]
  wire  _T_1687 = _T_1684 & _T_1686; // @[tlb.scala 50:46]
  wire [31:0] _T_1689 = {{16'd0}, tlb_entries_pagemask__T_1557_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1690 = ~_T_1689; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1415 = {{13'd0}, tlb_entries_vpn__T_1557_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1691 = _GEN_1415 & _T_1690; // @[tlb.scala 50:19]
  wire [31:0] _T_1693 = _GEN_1394 & _T_1690; // @[tlb.scala 50:37]
  wire  _T_1694 = _T_1691 == _T_1693; // @[tlb.scala 50:28]
  wire  _T_1695 = tlb_entries_asid__T_1557_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1696 = tlb_entries_g__T_1557_data | _T_1695; // @[tlb.scala 51:17]
  wire  _T_1697 = _T_1694 & _T_1696; // @[tlb.scala 50:46]
  wire [31:0] _T_1699 = {{16'd0}, tlb_entries_pagemask__T_1558_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1700 = ~_T_1699; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1417 = {{13'd0}, tlb_entries_vpn__T_1558_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1701 = _GEN_1417 & _T_1700; // @[tlb.scala 50:19]
  wire [31:0] _T_1703 = _GEN_1394 & _T_1700; // @[tlb.scala 50:37]
  wire  _T_1704 = _T_1701 == _T_1703; // @[tlb.scala 50:28]
  wire  _T_1705 = tlb_entries_asid__T_1558_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1706 = tlb_entries_g__T_1558_data | _T_1705; // @[tlb.scala 51:17]
  wire  _T_1707 = _T_1704 & _T_1706; // @[tlb.scala 50:46]
  wire [31:0] _T_1709 = {{16'd0}, tlb_entries_pagemask__T_1559_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1710 = ~_T_1709; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1419 = {{13'd0}, tlb_entries_vpn__T_1559_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1711 = _GEN_1419 & _T_1710; // @[tlb.scala 50:19]
  wire [31:0] _T_1713 = _GEN_1394 & _T_1710; // @[tlb.scala 50:37]
  wire  _T_1714 = _T_1711 == _T_1713; // @[tlb.scala 50:28]
  wire  _T_1715 = tlb_entries_asid__T_1559_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1716 = tlb_entries_g__T_1559_data | _T_1715; // @[tlb.scala 51:17]
  wire  _T_1717 = _T_1714 & _T_1716; // @[tlb.scala 50:46]
  wire [31:0] _T_1719 = {{16'd0}, tlb_entries_pagemask__T_1560_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1720 = ~_T_1719; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1421 = {{13'd0}, tlb_entries_vpn__T_1560_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1721 = _GEN_1421 & _T_1720; // @[tlb.scala 50:19]
  wire [31:0] _T_1723 = _GEN_1394 & _T_1720; // @[tlb.scala 50:37]
  wire  _T_1724 = _T_1721 == _T_1723; // @[tlb.scala 50:28]
  wire  _T_1725 = tlb_entries_asid__T_1560_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1726 = tlb_entries_g__T_1560_data | _T_1725; // @[tlb.scala 51:17]
  wire  _T_1727 = _T_1724 & _T_1726; // @[tlb.scala 50:46]
  wire [31:0] _T_1729 = {{16'd0}, tlb_entries_pagemask__T_1561_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1730 = ~_T_1729; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1423 = {{13'd0}, tlb_entries_vpn__T_1561_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1731 = _GEN_1423 & _T_1730; // @[tlb.scala 50:19]
  wire [31:0] _T_1733 = _GEN_1394 & _T_1730; // @[tlb.scala 50:37]
  wire  _T_1734 = _T_1731 == _T_1733; // @[tlb.scala 50:28]
  wire  _T_1735 = tlb_entries_asid__T_1561_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1736 = tlb_entries_g__T_1561_data | _T_1735; // @[tlb.scala 51:17]
  wire  _T_1737 = _T_1734 & _T_1736; // @[tlb.scala 50:46]
  wire [31:0] _T_1739 = {{16'd0}, tlb_entries_pagemask__T_1562_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1740 = ~_T_1739; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1425 = {{13'd0}, tlb_entries_vpn__T_1562_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1741 = _GEN_1425 & _T_1740; // @[tlb.scala 50:19]
  wire [31:0] _T_1743 = _GEN_1394 & _T_1740; // @[tlb.scala 50:37]
  wire  _T_1744 = _T_1741 == _T_1743; // @[tlb.scala 50:28]
  wire  _T_1745 = tlb_entries_asid__T_1562_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1746 = tlb_entries_g__T_1562_data | _T_1745; // @[tlb.scala 51:17]
  wire  _T_1747 = _T_1744 & _T_1746; // @[tlb.scala 50:46]
  wire [31:0] _T_1749 = {{16'd0}, tlb_entries_pagemask__T_1563_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1750 = ~_T_1749; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1427 = {{13'd0}, tlb_entries_vpn__T_1563_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1751 = _GEN_1427 & _T_1750; // @[tlb.scala 50:19]
  wire [31:0] _T_1753 = _GEN_1394 & _T_1750; // @[tlb.scala 50:37]
  wire  _T_1754 = _T_1751 == _T_1753; // @[tlb.scala 50:28]
  wire  _T_1755 = tlb_entries_asid__T_1563_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1756 = tlb_entries_g__T_1563_data | _T_1755; // @[tlb.scala 51:17]
  wire  _T_1757 = _T_1754 & _T_1756; // @[tlb.scala 50:46]
  wire [31:0] _T_1759 = {{16'd0}, tlb_entries_pagemask__T_1564_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1760 = ~_T_1759; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1429 = {{13'd0}, tlb_entries_vpn__T_1564_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1761 = _GEN_1429 & _T_1760; // @[tlb.scala 50:19]
  wire [31:0] _T_1763 = _GEN_1394 & _T_1760; // @[tlb.scala 50:37]
  wire  _T_1764 = _T_1761 == _T_1763; // @[tlb.scala 50:28]
  wire  _T_1765 = tlb_entries_asid__T_1564_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1766 = tlb_entries_g__T_1564_data | _T_1765; // @[tlb.scala 51:17]
  wire  _T_1767 = _T_1764 & _T_1766; // @[tlb.scala 50:46]
  wire [31:0] _T_1769 = {{16'd0}, tlb_entries_pagemask__T_1565_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1770 = ~_T_1769; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1431 = {{13'd0}, tlb_entries_vpn__T_1565_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1771 = _GEN_1431 & _T_1770; // @[tlb.scala 50:19]
  wire [31:0] _T_1773 = _GEN_1394 & _T_1770; // @[tlb.scala 50:37]
  wire  _T_1774 = _T_1771 == _T_1773; // @[tlb.scala 50:28]
  wire  _T_1775 = tlb_entries_asid__T_1565_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1776 = tlb_entries_g__T_1565_data | _T_1775; // @[tlb.scala 51:17]
  wire  _T_1777 = _T_1774 & _T_1776; // @[tlb.scala 50:46]
  wire [31:0] _T_1779 = {{16'd0}, tlb_entries_pagemask__T_1566_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1780 = ~_T_1779; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1433 = {{13'd0}, tlb_entries_vpn__T_1566_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1781 = _GEN_1433 & _T_1780; // @[tlb.scala 50:19]
  wire [31:0] _T_1783 = _GEN_1394 & _T_1780; // @[tlb.scala 50:37]
  wire  _T_1784 = _T_1781 == _T_1783; // @[tlb.scala 50:28]
  wire  _T_1785 = tlb_entries_asid__T_1566_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1786 = tlb_entries_g__T_1566_data | _T_1785; // @[tlb.scala 51:17]
  wire  _T_1787 = _T_1784 & _T_1786; // @[tlb.scala 50:46]
  wire [31:0] _T_1789 = {{16'd0}, tlb_entries_pagemask__T_1567_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1790 = ~_T_1789; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1435 = {{13'd0}, tlb_entries_vpn__T_1567_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1791 = _GEN_1435 & _T_1790; // @[tlb.scala 50:19]
  wire [31:0] _T_1793 = _GEN_1394 & _T_1790; // @[tlb.scala 50:37]
  wire  _T_1794 = _T_1791 == _T_1793; // @[tlb.scala 50:28]
  wire  _T_1795 = tlb_entries_asid__T_1567_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1796 = tlb_entries_g__T_1567_data | _T_1795; // @[tlb.scala 51:17]
  wire  _T_1797 = _T_1794 & _T_1796; // @[tlb.scala 50:46]
  wire [31:0] _T_1799 = {{16'd0}, tlb_entries_pagemask__T_1568_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1800 = ~_T_1799; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1437 = {{13'd0}, tlb_entries_vpn__T_1568_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1801 = _GEN_1437 & _T_1800; // @[tlb.scala 50:19]
  wire [31:0] _T_1803 = _GEN_1394 & _T_1800; // @[tlb.scala 50:37]
  wire  _T_1804 = _T_1801 == _T_1803; // @[tlb.scala 50:28]
  wire  _T_1805 = tlb_entries_asid__T_1568_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1806 = tlb_entries_g__T_1568_data | _T_1805; // @[tlb.scala 51:17]
  wire  _T_1807 = _T_1804 & _T_1806; // @[tlb.scala 50:46]
  wire [31:0] _T_1809 = {{16'd0}, tlb_entries_pagemask__T_1569_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1810 = ~_T_1809; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1439 = {{13'd0}, tlb_entries_vpn__T_1569_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1811 = _GEN_1439 & _T_1810; // @[tlb.scala 50:19]
  wire [31:0] _T_1813 = _GEN_1394 & _T_1810; // @[tlb.scala 50:37]
  wire  _T_1814 = _T_1811 == _T_1813; // @[tlb.scala 50:28]
  wire  _T_1815 = tlb_entries_asid__T_1569_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1816 = tlb_entries_g__T_1569_data | _T_1815; // @[tlb.scala 51:17]
  wire  _T_1817 = _T_1814 & _T_1816; // @[tlb.scala 50:46]
  wire [31:0] _T_1819 = {{16'd0}, tlb_entries_pagemask__T_1570_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1820 = ~_T_1819; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1441 = {{13'd0}, tlb_entries_vpn__T_1570_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1821 = _GEN_1441 & _T_1820; // @[tlb.scala 50:19]
  wire [31:0] _T_1823 = _GEN_1394 & _T_1820; // @[tlb.scala 50:37]
  wire  _T_1824 = _T_1821 == _T_1823; // @[tlb.scala 50:28]
  wire  _T_1825 = tlb_entries_asid__T_1570_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1826 = tlb_entries_g__T_1570_data | _T_1825; // @[tlb.scala 51:17]
  wire  _T_1827 = _T_1824 & _T_1826; // @[tlb.scala 50:46]
  wire [31:0] _T_1829 = {{16'd0}, tlb_entries_pagemask__T_1571_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1830 = ~_T_1829; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1443 = {{13'd0}, tlb_entries_vpn__T_1571_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1831 = _GEN_1443 & _T_1830; // @[tlb.scala 50:19]
  wire [31:0] _T_1833 = _GEN_1394 & _T_1830; // @[tlb.scala 50:37]
  wire  _T_1834 = _T_1831 == _T_1833; // @[tlb.scala 50:28]
  wire  _T_1835 = tlb_entries_asid__T_1571_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1836 = tlb_entries_g__T_1571_data | _T_1835; // @[tlb.scala 51:17]
  wire  _T_1837 = _T_1834 & _T_1836; // @[tlb.scala 50:46]
  wire [31:0] _T_1839 = {{16'd0}, tlb_entries_pagemask__T_1572_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1840 = ~_T_1839; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1445 = {{13'd0}, tlb_entries_vpn__T_1572_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1841 = _GEN_1445 & _T_1840; // @[tlb.scala 50:19]
  wire [31:0] _T_1843 = _GEN_1394 & _T_1840; // @[tlb.scala 50:37]
  wire  _T_1844 = _T_1841 == _T_1843; // @[tlb.scala 50:28]
  wire  _T_1845 = tlb_entries_asid__T_1572_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1846 = tlb_entries_g__T_1572_data | _T_1845; // @[tlb.scala 51:17]
  wire  _T_1847 = _T_1844 & _T_1846; // @[tlb.scala 50:46]
  wire [31:0] _T_1849 = {{16'd0}, tlb_entries_pagemask__T_1573_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1850 = ~_T_1849; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1447 = {{13'd0}, tlb_entries_vpn__T_1573_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1851 = _GEN_1447 & _T_1850; // @[tlb.scala 50:19]
  wire [31:0] _T_1853 = _GEN_1394 & _T_1850; // @[tlb.scala 50:37]
  wire  _T_1854 = _T_1851 == _T_1853; // @[tlb.scala 50:28]
  wire  _T_1855 = tlb_entries_asid__T_1573_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1856 = tlb_entries_g__T_1573_data | _T_1855; // @[tlb.scala 51:17]
  wire  _T_1857 = _T_1854 & _T_1856; // @[tlb.scala 50:46]
  wire [31:0] _T_1859 = {{16'd0}, tlb_entries_pagemask__T_1574_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1860 = ~_T_1859; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1449 = {{13'd0}, tlb_entries_vpn__T_1574_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1861 = _GEN_1449 & _T_1860; // @[tlb.scala 50:19]
  wire [31:0] _T_1863 = _GEN_1394 & _T_1860; // @[tlb.scala 50:37]
  wire  _T_1864 = _T_1861 == _T_1863; // @[tlb.scala 50:28]
  wire  _T_1865 = tlb_entries_asid__T_1574_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1866 = tlb_entries_g__T_1574_data | _T_1865; // @[tlb.scala 51:17]
  wire  _T_1867 = _T_1864 & _T_1866; // @[tlb.scala 50:46]
  wire [31:0] _T_1869 = {{16'd0}, tlb_entries_pagemask__T_1575_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1870 = ~_T_1869; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1451 = {{13'd0}, tlb_entries_vpn__T_1575_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1871 = _GEN_1451 & _T_1870; // @[tlb.scala 50:19]
  wire [31:0] _T_1873 = _GEN_1394 & _T_1870; // @[tlb.scala 50:37]
  wire  _T_1874 = _T_1871 == _T_1873; // @[tlb.scala 50:28]
  wire  _T_1875 = tlb_entries_asid__T_1575_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1876 = tlb_entries_g__T_1575_data | _T_1875; // @[tlb.scala 51:17]
  wire  _T_1877 = _T_1874 & _T_1876; // @[tlb.scala 50:46]
  wire [31:0] _T_1879 = {{16'd0}, tlb_entries_pagemask__T_1576_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1880 = ~_T_1879; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1453 = {{13'd0}, tlb_entries_vpn__T_1576_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1881 = _GEN_1453 & _T_1880; // @[tlb.scala 50:19]
  wire [31:0] _T_1883 = _GEN_1394 & _T_1880; // @[tlb.scala 50:37]
  wire  _T_1884 = _T_1881 == _T_1883; // @[tlb.scala 50:28]
  wire  _T_1885 = tlb_entries_asid__T_1576_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1886 = tlb_entries_g__T_1576_data | _T_1885; // @[tlb.scala 51:17]
  wire  _T_1887 = _T_1884 & _T_1886; // @[tlb.scala 50:46]
  wire [31:0] _T_1889 = {{16'd0}, tlb_entries_pagemask__T_1577_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_1890 = ~_T_1889; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1455 = {{13'd0}, tlb_entries_vpn__T_1577_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_1891 = _GEN_1455 & _T_1890; // @[tlb.scala 50:19]
  wire [31:0] _T_1893 = _GEN_1394 & _T_1890; // @[tlb.scala 50:37]
  wire  _T_1894 = _T_1891 == _T_1893; // @[tlb.scala 50:28]
  wire  _T_1895 = tlb_entries_asid__T_1577_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_1896 = tlb_entries_g__T_1577_data | _T_1895; // @[tlb.scala 51:17]
  wire  _T_1897 = _T_1894 & _T_1896; // @[tlb.scala 50:46]
  wire [7:0] _T_1904 = {_T_1827,_T_1837,_T_1847,_T_1857,_T_1867,_T_1877,_T_1887,_T_1897}; // @[Cat.scala 29:58]
  wire [15:0] _T_1912 = {_T_1747,_T_1757,_T_1767,_T_1777,_T_1787,_T_1797,_T_1807,_T_1817,_T_1904}; // @[Cat.scala 29:58]
  wire [7:0] _T_1919 = {_T_1667,_T_1677,_T_1687,_T_1697,_T_1707,_T_1717,_T_1727,_T_1737}; // @[Cat.scala 29:58]
  wire [31:0] _T_1928 = {_T_1587,_T_1597,_T_1607,_T_1617,_T_1627,_T_1637,_T_1647,_T_1657,_T_1919,_T_1912}; // @[Cat.scala 29:58]
  wire [31:0] _T_1932 = {{16'd0}, _T_1928[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1934 = {_T_1928[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1936 = _T_1934 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1937 = _T_1932 | _T_1936; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1457 = {{8'd0}, _T_1937[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1942 = _GEN_1457 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1944 = {_T_1937[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1946 = _T_1944 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1947 = _T_1942 | _T_1946; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1458 = {{4'd0}, _T_1947[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1952 = _GEN_1458 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1954 = {_T_1947[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1956 = _T_1954 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1957 = _T_1952 | _T_1956; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1459 = {{2'd0}, _T_1957[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1962 = _GEN_1459 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1964 = {_T_1957[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1966 = _T_1964 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1967 = _T_1962 | _T_1966; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1460 = {{1'd0}, _T_1967[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1972 = _GEN_1460 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_1974 = {_T_1967[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_1976 = _T_1974 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_1977 = _T_1972 | _T_1976; // @[Bitwise.scala 103:39]
  wire  _T_1978 = _T_1977 != 32'h0; // @[tlb.scala 83:25]
  wire  _T_1979 = ~_T_1978; // @[tlb.scala 83:16]
  wire [31:0] _T_1983 = _T_1579 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_1984 = {_T_1983, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _GEN_1461 = {{12'd0}, _T_1544_vaddr}; // @[tlb.scala 55:24]
  wire [43:0] _T_1985 = _GEN_1461 & _T_1984; // @[tlb.scala 55:24]
  wire  _T_1986 = _T_1985 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_1987_pfn = _T_1986 ? tlb_entries_p1_pfn__T_1546_data : tlb_entries_p0_pfn__T_1546_data; // @[tlb.scala 56:19]
  wire  _T_1987_d = _T_1986 ? tlb_entries_p1_d__T_1546_data : tlb_entries_p0_d__T_1546_data; // @[tlb.scala 56:19]
  wire  _T_1987_v = _T_1986 ? tlb_entries_p1_v__T_1546_data : tlb_entries_p0_v__T_1546_data; // @[tlb.scala 56:19]
  wire  _T_1988 = ~_T_1544_func; // @[tlb.scala 57:28]
  wire [4:0] _T_1989 = _T_1988 ? 5'h2 : 5'h3; // @[tlb.scala 57:21]
  wire  _T_1992 = ~_T_1987_v; // @[tlb.scala 59:18]
  wire  _T_1993 = ~_T_1987_d; // @[tlb.scala 63:25]
  wire  _T_1995 = _T_1993 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1462 = {{8'd0}, _T_1987_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_1997 = _GEN_1462 & _T_1580; // @[tlb.scala 68:32]
  wire [43:0] _T_1998 = {_T_1997, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2003 = _T_1984 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2004 = _GEN_1461 & _T_2003; // @[tlb.scala 69:27]
  wire [43:0] _T_2005 = _T_1998 | _T_2004; // @[tlb.scala 70:29]
  wire [4:0] _GEN_202 = _T_1995 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_203 = _T_1995 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_204 = _T_1995 ? 44'h0 : _T_2005; // @[tlb.scala 63:53]
  wire [4:0] _GEN_205 = _T_1992 ? 5'h8 : _GEN_202; // @[tlb.scala 59:27]
  wire [4:0] _GEN_206 = _T_1992 ? _T_1989 : _GEN_203; // @[tlb.scala 59:27]
  wire [43:0] _GEN_207 = _T_1992 ? 44'h0 : _GEN_204; // @[tlb.scala 59:27]
  wire [31:0] _T_2009 = _T_1589 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2010 = {_T_2009, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2011 = _GEN_1461 & _T_2010; // @[tlb.scala 55:24]
  wire  _T_2012 = _T_2011 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2013_pfn = _T_2012 ? tlb_entries_p1_pfn__T_1547_data : tlb_entries_p0_pfn__T_1547_data; // @[tlb.scala 56:19]
  wire  _T_2013_d = _T_2012 ? tlb_entries_p1_d__T_1547_data : tlb_entries_p0_d__T_1547_data; // @[tlb.scala 56:19]
  wire  _T_2013_v = _T_2012 ? tlb_entries_p1_v__T_1547_data : tlb_entries_p0_v__T_1547_data; // @[tlb.scala 56:19]
  wire  _T_2018 = ~_T_2013_v; // @[tlb.scala 59:18]
  wire  _T_2019 = ~_T_2013_d; // @[tlb.scala 63:25]
  wire  _T_2021 = _T_2019 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1465 = {{8'd0}, _T_2013_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2023 = _GEN_1465 & _T_1590; // @[tlb.scala 68:32]
  wire [43:0] _T_2024 = {_T_2023, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2029 = _T_2010 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2030 = _GEN_1461 & _T_2029; // @[tlb.scala 69:27]
  wire [43:0] _T_2031 = _T_2024 | _T_2030; // @[tlb.scala 70:29]
  wire [4:0] _GEN_208 = _T_2021 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_209 = _T_2021 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_210 = _T_2021 ? 44'h0 : _T_2031; // @[tlb.scala 63:53]
  wire [4:0] _GEN_211 = _T_2018 ? 5'h8 : _GEN_208; // @[tlb.scala 59:27]
  wire [4:0] _GEN_212 = _T_2018 ? _T_1989 : _GEN_209; // @[tlb.scala 59:27]
  wire [43:0] _GEN_213 = _T_2018 ? 44'h0 : _GEN_210; // @[tlb.scala 59:27]
  wire [31:0] _T_2035 = _T_1599 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2036 = {_T_2035, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2037 = _GEN_1461 & _T_2036; // @[tlb.scala 55:24]
  wire  _T_2038 = _T_2037 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2039_pfn = _T_2038 ? tlb_entries_p1_pfn__T_1548_data : tlb_entries_p0_pfn__T_1548_data; // @[tlb.scala 56:19]
  wire  _T_2039_d = _T_2038 ? tlb_entries_p1_d__T_1548_data : tlb_entries_p0_d__T_1548_data; // @[tlb.scala 56:19]
  wire  _T_2039_v = _T_2038 ? tlb_entries_p1_v__T_1548_data : tlb_entries_p0_v__T_1548_data; // @[tlb.scala 56:19]
  wire  _T_2044 = ~_T_2039_v; // @[tlb.scala 59:18]
  wire  _T_2045 = ~_T_2039_d; // @[tlb.scala 63:25]
  wire  _T_2047 = _T_2045 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1468 = {{8'd0}, _T_2039_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2049 = _GEN_1468 & _T_1600; // @[tlb.scala 68:32]
  wire [43:0] _T_2050 = {_T_2049, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2055 = _T_2036 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2056 = _GEN_1461 & _T_2055; // @[tlb.scala 69:27]
  wire [43:0] _T_2057 = _T_2050 | _T_2056; // @[tlb.scala 70:29]
  wire [4:0] _GEN_214 = _T_2047 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_215 = _T_2047 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_216 = _T_2047 ? 44'h0 : _T_2057; // @[tlb.scala 63:53]
  wire [4:0] _GEN_217 = _T_2044 ? 5'h8 : _GEN_214; // @[tlb.scala 59:27]
  wire [4:0] _GEN_218 = _T_2044 ? _T_1989 : _GEN_215; // @[tlb.scala 59:27]
  wire [43:0] _GEN_219 = _T_2044 ? 44'h0 : _GEN_216; // @[tlb.scala 59:27]
  wire [31:0] _T_2061 = _T_1609 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2062 = {_T_2061, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2063 = _GEN_1461 & _T_2062; // @[tlb.scala 55:24]
  wire  _T_2064 = _T_2063 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2065_pfn = _T_2064 ? tlb_entries_p1_pfn__T_1549_data : tlb_entries_p0_pfn__T_1549_data; // @[tlb.scala 56:19]
  wire  _T_2065_d = _T_2064 ? tlb_entries_p1_d__T_1549_data : tlb_entries_p0_d__T_1549_data; // @[tlb.scala 56:19]
  wire  _T_2065_v = _T_2064 ? tlb_entries_p1_v__T_1549_data : tlb_entries_p0_v__T_1549_data; // @[tlb.scala 56:19]
  wire  _T_2070 = ~_T_2065_v; // @[tlb.scala 59:18]
  wire  _T_2071 = ~_T_2065_d; // @[tlb.scala 63:25]
  wire  _T_2073 = _T_2071 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1471 = {{8'd0}, _T_2065_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2075 = _GEN_1471 & _T_1610; // @[tlb.scala 68:32]
  wire [43:0] _T_2076 = {_T_2075, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2081 = _T_2062 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2082 = _GEN_1461 & _T_2081; // @[tlb.scala 69:27]
  wire [43:0] _T_2083 = _T_2076 | _T_2082; // @[tlb.scala 70:29]
  wire [4:0] _GEN_220 = _T_2073 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_221 = _T_2073 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_222 = _T_2073 ? 44'h0 : _T_2083; // @[tlb.scala 63:53]
  wire [4:0] _GEN_223 = _T_2070 ? 5'h8 : _GEN_220; // @[tlb.scala 59:27]
  wire [4:0] _GEN_224 = _T_2070 ? _T_1989 : _GEN_221; // @[tlb.scala 59:27]
  wire [43:0] _GEN_225 = _T_2070 ? 44'h0 : _GEN_222; // @[tlb.scala 59:27]
  wire [31:0] _T_2087 = _T_1619 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2088 = {_T_2087, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2089 = _GEN_1461 & _T_2088; // @[tlb.scala 55:24]
  wire  _T_2090 = _T_2089 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2091_pfn = _T_2090 ? tlb_entries_p1_pfn__T_1550_data : tlb_entries_p0_pfn__T_1550_data; // @[tlb.scala 56:19]
  wire  _T_2091_d = _T_2090 ? tlb_entries_p1_d__T_1550_data : tlb_entries_p0_d__T_1550_data; // @[tlb.scala 56:19]
  wire  _T_2091_v = _T_2090 ? tlb_entries_p1_v__T_1550_data : tlb_entries_p0_v__T_1550_data; // @[tlb.scala 56:19]
  wire  _T_2096 = ~_T_2091_v; // @[tlb.scala 59:18]
  wire  _T_2097 = ~_T_2091_d; // @[tlb.scala 63:25]
  wire  _T_2099 = _T_2097 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1474 = {{8'd0}, _T_2091_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2101 = _GEN_1474 & _T_1620; // @[tlb.scala 68:32]
  wire [43:0] _T_2102 = {_T_2101, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2107 = _T_2088 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2108 = _GEN_1461 & _T_2107; // @[tlb.scala 69:27]
  wire [43:0] _T_2109 = _T_2102 | _T_2108; // @[tlb.scala 70:29]
  wire [4:0] _GEN_226 = _T_2099 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_227 = _T_2099 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_228 = _T_2099 ? 44'h0 : _T_2109; // @[tlb.scala 63:53]
  wire [4:0] _GEN_229 = _T_2096 ? 5'h8 : _GEN_226; // @[tlb.scala 59:27]
  wire [4:0] _GEN_230 = _T_2096 ? _T_1989 : _GEN_227; // @[tlb.scala 59:27]
  wire [43:0] _GEN_231 = _T_2096 ? 44'h0 : _GEN_228; // @[tlb.scala 59:27]
  wire [31:0] _T_2113 = _T_1629 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2114 = {_T_2113, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2115 = _GEN_1461 & _T_2114; // @[tlb.scala 55:24]
  wire  _T_2116 = _T_2115 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2117_pfn = _T_2116 ? tlb_entries_p1_pfn__T_1551_data : tlb_entries_p0_pfn__T_1551_data; // @[tlb.scala 56:19]
  wire  _T_2117_d = _T_2116 ? tlb_entries_p1_d__T_1551_data : tlb_entries_p0_d__T_1551_data; // @[tlb.scala 56:19]
  wire  _T_2117_v = _T_2116 ? tlb_entries_p1_v__T_1551_data : tlb_entries_p0_v__T_1551_data; // @[tlb.scala 56:19]
  wire  _T_2122 = ~_T_2117_v; // @[tlb.scala 59:18]
  wire  _T_2123 = ~_T_2117_d; // @[tlb.scala 63:25]
  wire  _T_2125 = _T_2123 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1477 = {{8'd0}, _T_2117_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2127 = _GEN_1477 & _T_1630; // @[tlb.scala 68:32]
  wire [43:0] _T_2128 = {_T_2127, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2133 = _T_2114 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2134 = _GEN_1461 & _T_2133; // @[tlb.scala 69:27]
  wire [43:0] _T_2135 = _T_2128 | _T_2134; // @[tlb.scala 70:29]
  wire [4:0] _GEN_232 = _T_2125 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_233 = _T_2125 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_234 = _T_2125 ? 44'h0 : _T_2135; // @[tlb.scala 63:53]
  wire [4:0] _GEN_235 = _T_2122 ? 5'h8 : _GEN_232; // @[tlb.scala 59:27]
  wire [4:0] _GEN_236 = _T_2122 ? _T_1989 : _GEN_233; // @[tlb.scala 59:27]
  wire [43:0] _GEN_237 = _T_2122 ? 44'h0 : _GEN_234; // @[tlb.scala 59:27]
  wire [31:0] _T_2139 = _T_1639 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2140 = {_T_2139, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2141 = _GEN_1461 & _T_2140; // @[tlb.scala 55:24]
  wire  _T_2142 = _T_2141 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2143_pfn = _T_2142 ? tlb_entries_p1_pfn__T_1552_data : tlb_entries_p0_pfn__T_1552_data; // @[tlb.scala 56:19]
  wire  _T_2143_d = _T_2142 ? tlb_entries_p1_d__T_1552_data : tlb_entries_p0_d__T_1552_data; // @[tlb.scala 56:19]
  wire  _T_2143_v = _T_2142 ? tlb_entries_p1_v__T_1552_data : tlb_entries_p0_v__T_1552_data; // @[tlb.scala 56:19]
  wire  _T_2148 = ~_T_2143_v; // @[tlb.scala 59:18]
  wire  _T_2149 = ~_T_2143_d; // @[tlb.scala 63:25]
  wire  _T_2151 = _T_2149 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1480 = {{8'd0}, _T_2143_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2153 = _GEN_1480 & _T_1640; // @[tlb.scala 68:32]
  wire [43:0] _T_2154 = {_T_2153, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2159 = _T_2140 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2160 = _GEN_1461 & _T_2159; // @[tlb.scala 69:27]
  wire [43:0] _T_2161 = _T_2154 | _T_2160; // @[tlb.scala 70:29]
  wire [4:0] _GEN_238 = _T_2151 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_239 = _T_2151 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_240 = _T_2151 ? 44'h0 : _T_2161; // @[tlb.scala 63:53]
  wire [4:0] _GEN_241 = _T_2148 ? 5'h8 : _GEN_238; // @[tlb.scala 59:27]
  wire [4:0] _GEN_242 = _T_2148 ? _T_1989 : _GEN_239; // @[tlb.scala 59:27]
  wire [43:0] _GEN_243 = _T_2148 ? 44'h0 : _GEN_240; // @[tlb.scala 59:27]
  wire [31:0] _T_2165 = _T_1649 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2166 = {_T_2165, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2167 = _GEN_1461 & _T_2166; // @[tlb.scala 55:24]
  wire  _T_2168 = _T_2167 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2169_pfn = _T_2168 ? tlb_entries_p1_pfn__T_1553_data : tlb_entries_p0_pfn__T_1553_data; // @[tlb.scala 56:19]
  wire  _T_2169_d = _T_2168 ? tlb_entries_p1_d__T_1553_data : tlb_entries_p0_d__T_1553_data; // @[tlb.scala 56:19]
  wire  _T_2169_v = _T_2168 ? tlb_entries_p1_v__T_1553_data : tlb_entries_p0_v__T_1553_data; // @[tlb.scala 56:19]
  wire  _T_2174 = ~_T_2169_v; // @[tlb.scala 59:18]
  wire  _T_2175 = ~_T_2169_d; // @[tlb.scala 63:25]
  wire  _T_2177 = _T_2175 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1483 = {{8'd0}, _T_2169_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2179 = _GEN_1483 & _T_1650; // @[tlb.scala 68:32]
  wire [43:0] _T_2180 = {_T_2179, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2185 = _T_2166 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2186 = _GEN_1461 & _T_2185; // @[tlb.scala 69:27]
  wire [43:0] _T_2187 = _T_2180 | _T_2186; // @[tlb.scala 70:29]
  wire [4:0] _GEN_244 = _T_2177 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_245 = _T_2177 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_246 = _T_2177 ? 44'h0 : _T_2187; // @[tlb.scala 63:53]
  wire [4:0] _GEN_247 = _T_2174 ? 5'h8 : _GEN_244; // @[tlb.scala 59:27]
  wire [4:0] _GEN_248 = _T_2174 ? _T_1989 : _GEN_245; // @[tlb.scala 59:27]
  wire [43:0] _GEN_249 = _T_2174 ? 44'h0 : _GEN_246; // @[tlb.scala 59:27]
  wire [31:0] _T_2191 = _T_1659 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2192 = {_T_2191, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2193 = _GEN_1461 & _T_2192; // @[tlb.scala 55:24]
  wire  _T_2194 = _T_2193 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2195_pfn = _T_2194 ? tlb_entries_p1_pfn__T_1554_data : tlb_entries_p0_pfn__T_1554_data; // @[tlb.scala 56:19]
  wire  _T_2195_d = _T_2194 ? tlb_entries_p1_d__T_1554_data : tlb_entries_p0_d__T_1554_data; // @[tlb.scala 56:19]
  wire  _T_2195_v = _T_2194 ? tlb_entries_p1_v__T_1554_data : tlb_entries_p0_v__T_1554_data; // @[tlb.scala 56:19]
  wire  _T_2200 = ~_T_2195_v; // @[tlb.scala 59:18]
  wire  _T_2201 = ~_T_2195_d; // @[tlb.scala 63:25]
  wire  _T_2203 = _T_2201 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1486 = {{8'd0}, _T_2195_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2205 = _GEN_1486 & _T_1660; // @[tlb.scala 68:32]
  wire [43:0] _T_2206 = {_T_2205, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2211 = _T_2192 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2212 = _GEN_1461 & _T_2211; // @[tlb.scala 69:27]
  wire [43:0] _T_2213 = _T_2206 | _T_2212; // @[tlb.scala 70:29]
  wire [4:0] _GEN_250 = _T_2203 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_251 = _T_2203 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_252 = _T_2203 ? 44'h0 : _T_2213; // @[tlb.scala 63:53]
  wire [4:0] _GEN_253 = _T_2200 ? 5'h8 : _GEN_250; // @[tlb.scala 59:27]
  wire [4:0] _GEN_254 = _T_2200 ? _T_1989 : _GEN_251; // @[tlb.scala 59:27]
  wire [43:0] _GEN_255 = _T_2200 ? 44'h0 : _GEN_252; // @[tlb.scala 59:27]
  wire [31:0] _T_2217 = _T_1669 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2218 = {_T_2217, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2219 = _GEN_1461 & _T_2218; // @[tlb.scala 55:24]
  wire  _T_2220 = _T_2219 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2221_pfn = _T_2220 ? tlb_entries_p1_pfn__T_1555_data : tlb_entries_p0_pfn__T_1555_data; // @[tlb.scala 56:19]
  wire  _T_2221_d = _T_2220 ? tlb_entries_p1_d__T_1555_data : tlb_entries_p0_d__T_1555_data; // @[tlb.scala 56:19]
  wire  _T_2221_v = _T_2220 ? tlb_entries_p1_v__T_1555_data : tlb_entries_p0_v__T_1555_data; // @[tlb.scala 56:19]
  wire  _T_2226 = ~_T_2221_v; // @[tlb.scala 59:18]
  wire  _T_2227 = ~_T_2221_d; // @[tlb.scala 63:25]
  wire  _T_2229 = _T_2227 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1489 = {{8'd0}, _T_2221_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2231 = _GEN_1489 & _T_1670; // @[tlb.scala 68:32]
  wire [43:0] _T_2232 = {_T_2231, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2237 = _T_2218 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2238 = _GEN_1461 & _T_2237; // @[tlb.scala 69:27]
  wire [43:0] _T_2239 = _T_2232 | _T_2238; // @[tlb.scala 70:29]
  wire [4:0] _GEN_256 = _T_2229 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_257 = _T_2229 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_258 = _T_2229 ? 44'h0 : _T_2239; // @[tlb.scala 63:53]
  wire [4:0] _GEN_259 = _T_2226 ? 5'h8 : _GEN_256; // @[tlb.scala 59:27]
  wire [4:0] _GEN_260 = _T_2226 ? _T_1989 : _GEN_257; // @[tlb.scala 59:27]
  wire [43:0] _GEN_261 = _T_2226 ? 44'h0 : _GEN_258; // @[tlb.scala 59:27]
  wire [31:0] _T_2243 = _T_1679 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2244 = {_T_2243, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2245 = _GEN_1461 & _T_2244; // @[tlb.scala 55:24]
  wire  _T_2246 = _T_2245 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2247_pfn = _T_2246 ? tlb_entries_p1_pfn__T_1556_data : tlb_entries_p0_pfn__T_1556_data; // @[tlb.scala 56:19]
  wire  _T_2247_d = _T_2246 ? tlb_entries_p1_d__T_1556_data : tlb_entries_p0_d__T_1556_data; // @[tlb.scala 56:19]
  wire  _T_2247_v = _T_2246 ? tlb_entries_p1_v__T_1556_data : tlb_entries_p0_v__T_1556_data; // @[tlb.scala 56:19]
  wire  _T_2252 = ~_T_2247_v; // @[tlb.scala 59:18]
  wire  _T_2253 = ~_T_2247_d; // @[tlb.scala 63:25]
  wire  _T_2255 = _T_2253 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1492 = {{8'd0}, _T_2247_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2257 = _GEN_1492 & _T_1680; // @[tlb.scala 68:32]
  wire [43:0] _T_2258 = {_T_2257, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2263 = _T_2244 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2264 = _GEN_1461 & _T_2263; // @[tlb.scala 69:27]
  wire [43:0] _T_2265 = _T_2258 | _T_2264; // @[tlb.scala 70:29]
  wire [4:0] _GEN_262 = _T_2255 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_263 = _T_2255 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_264 = _T_2255 ? 44'h0 : _T_2265; // @[tlb.scala 63:53]
  wire [4:0] _GEN_265 = _T_2252 ? 5'h8 : _GEN_262; // @[tlb.scala 59:27]
  wire [4:0] _GEN_266 = _T_2252 ? _T_1989 : _GEN_263; // @[tlb.scala 59:27]
  wire [43:0] _GEN_267 = _T_2252 ? 44'h0 : _GEN_264; // @[tlb.scala 59:27]
  wire [31:0] _T_2269 = _T_1689 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2270 = {_T_2269, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2271 = _GEN_1461 & _T_2270; // @[tlb.scala 55:24]
  wire  _T_2272 = _T_2271 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2273_pfn = _T_2272 ? tlb_entries_p1_pfn__T_1557_data : tlb_entries_p0_pfn__T_1557_data; // @[tlb.scala 56:19]
  wire  _T_2273_d = _T_2272 ? tlb_entries_p1_d__T_1557_data : tlb_entries_p0_d__T_1557_data; // @[tlb.scala 56:19]
  wire  _T_2273_v = _T_2272 ? tlb_entries_p1_v__T_1557_data : tlb_entries_p0_v__T_1557_data; // @[tlb.scala 56:19]
  wire  _T_2278 = ~_T_2273_v; // @[tlb.scala 59:18]
  wire  _T_2279 = ~_T_2273_d; // @[tlb.scala 63:25]
  wire  _T_2281 = _T_2279 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1495 = {{8'd0}, _T_2273_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2283 = _GEN_1495 & _T_1690; // @[tlb.scala 68:32]
  wire [43:0] _T_2284 = {_T_2283, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2289 = _T_2270 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2290 = _GEN_1461 & _T_2289; // @[tlb.scala 69:27]
  wire [43:0] _T_2291 = _T_2284 | _T_2290; // @[tlb.scala 70:29]
  wire [4:0] _GEN_268 = _T_2281 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_269 = _T_2281 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_270 = _T_2281 ? 44'h0 : _T_2291; // @[tlb.scala 63:53]
  wire [4:0] _GEN_271 = _T_2278 ? 5'h8 : _GEN_268; // @[tlb.scala 59:27]
  wire [4:0] _GEN_272 = _T_2278 ? _T_1989 : _GEN_269; // @[tlb.scala 59:27]
  wire [43:0] _GEN_273 = _T_2278 ? 44'h0 : _GEN_270; // @[tlb.scala 59:27]
  wire [31:0] _T_2295 = _T_1699 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2296 = {_T_2295, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2297 = _GEN_1461 & _T_2296; // @[tlb.scala 55:24]
  wire  _T_2298 = _T_2297 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2299_pfn = _T_2298 ? tlb_entries_p1_pfn__T_1558_data : tlb_entries_p0_pfn__T_1558_data; // @[tlb.scala 56:19]
  wire  _T_2299_d = _T_2298 ? tlb_entries_p1_d__T_1558_data : tlb_entries_p0_d__T_1558_data; // @[tlb.scala 56:19]
  wire  _T_2299_v = _T_2298 ? tlb_entries_p1_v__T_1558_data : tlb_entries_p0_v__T_1558_data; // @[tlb.scala 56:19]
  wire  _T_2304 = ~_T_2299_v; // @[tlb.scala 59:18]
  wire  _T_2305 = ~_T_2299_d; // @[tlb.scala 63:25]
  wire  _T_2307 = _T_2305 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1498 = {{8'd0}, _T_2299_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2309 = _GEN_1498 & _T_1700; // @[tlb.scala 68:32]
  wire [43:0] _T_2310 = {_T_2309, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2315 = _T_2296 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2316 = _GEN_1461 & _T_2315; // @[tlb.scala 69:27]
  wire [43:0] _T_2317 = _T_2310 | _T_2316; // @[tlb.scala 70:29]
  wire [4:0] _GEN_274 = _T_2307 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_275 = _T_2307 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_276 = _T_2307 ? 44'h0 : _T_2317; // @[tlb.scala 63:53]
  wire [4:0] _GEN_277 = _T_2304 ? 5'h8 : _GEN_274; // @[tlb.scala 59:27]
  wire [4:0] _GEN_278 = _T_2304 ? _T_1989 : _GEN_275; // @[tlb.scala 59:27]
  wire [43:0] _GEN_279 = _T_2304 ? 44'h0 : _GEN_276; // @[tlb.scala 59:27]
  wire [31:0] _T_2321 = _T_1709 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2322 = {_T_2321, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2323 = _GEN_1461 & _T_2322; // @[tlb.scala 55:24]
  wire  _T_2324 = _T_2323 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2325_pfn = _T_2324 ? tlb_entries_p1_pfn__T_1559_data : tlb_entries_p0_pfn__T_1559_data; // @[tlb.scala 56:19]
  wire  _T_2325_d = _T_2324 ? tlb_entries_p1_d__T_1559_data : tlb_entries_p0_d__T_1559_data; // @[tlb.scala 56:19]
  wire  _T_2325_v = _T_2324 ? tlb_entries_p1_v__T_1559_data : tlb_entries_p0_v__T_1559_data; // @[tlb.scala 56:19]
  wire  _T_2330 = ~_T_2325_v; // @[tlb.scala 59:18]
  wire  _T_2331 = ~_T_2325_d; // @[tlb.scala 63:25]
  wire  _T_2333 = _T_2331 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1501 = {{8'd0}, _T_2325_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2335 = _GEN_1501 & _T_1710; // @[tlb.scala 68:32]
  wire [43:0] _T_2336 = {_T_2335, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2341 = _T_2322 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2342 = _GEN_1461 & _T_2341; // @[tlb.scala 69:27]
  wire [43:0] _T_2343 = _T_2336 | _T_2342; // @[tlb.scala 70:29]
  wire [4:0] _GEN_280 = _T_2333 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_281 = _T_2333 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_282 = _T_2333 ? 44'h0 : _T_2343; // @[tlb.scala 63:53]
  wire [4:0] _GEN_283 = _T_2330 ? 5'h8 : _GEN_280; // @[tlb.scala 59:27]
  wire [4:0] _GEN_284 = _T_2330 ? _T_1989 : _GEN_281; // @[tlb.scala 59:27]
  wire [43:0] _GEN_285 = _T_2330 ? 44'h0 : _GEN_282; // @[tlb.scala 59:27]
  wire [31:0] _T_2347 = _T_1719 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2348 = {_T_2347, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2349 = _GEN_1461 & _T_2348; // @[tlb.scala 55:24]
  wire  _T_2350 = _T_2349 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2351_pfn = _T_2350 ? tlb_entries_p1_pfn__T_1560_data : tlb_entries_p0_pfn__T_1560_data; // @[tlb.scala 56:19]
  wire  _T_2351_d = _T_2350 ? tlb_entries_p1_d__T_1560_data : tlb_entries_p0_d__T_1560_data; // @[tlb.scala 56:19]
  wire  _T_2351_v = _T_2350 ? tlb_entries_p1_v__T_1560_data : tlb_entries_p0_v__T_1560_data; // @[tlb.scala 56:19]
  wire  _T_2356 = ~_T_2351_v; // @[tlb.scala 59:18]
  wire  _T_2357 = ~_T_2351_d; // @[tlb.scala 63:25]
  wire  _T_2359 = _T_2357 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1504 = {{8'd0}, _T_2351_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2361 = _GEN_1504 & _T_1720; // @[tlb.scala 68:32]
  wire [43:0] _T_2362 = {_T_2361, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2367 = _T_2348 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2368 = _GEN_1461 & _T_2367; // @[tlb.scala 69:27]
  wire [43:0] _T_2369 = _T_2362 | _T_2368; // @[tlb.scala 70:29]
  wire [4:0] _GEN_286 = _T_2359 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_287 = _T_2359 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_288 = _T_2359 ? 44'h0 : _T_2369; // @[tlb.scala 63:53]
  wire [4:0] _GEN_289 = _T_2356 ? 5'h8 : _GEN_286; // @[tlb.scala 59:27]
  wire [4:0] _GEN_290 = _T_2356 ? _T_1989 : _GEN_287; // @[tlb.scala 59:27]
  wire [43:0] _GEN_291 = _T_2356 ? 44'h0 : _GEN_288; // @[tlb.scala 59:27]
  wire [31:0] _T_2373 = _T_1729 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2374 = {_T_2373, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2375 = _GEN_1461 & _T_2374; // @[tlb.scala 55:24]
  wire  _T_2376 = _T_2375 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2377_pfn = _T_2376 ? tlb_entries_p1_pfn__T_1561_data : tlb_entries_p0_pfn__T_1561_data; // @[tlb.scala 56:19]
  wire  _T_2377_d = _T_2376 ? tlb_entries_p1_d__T_1561_data : tlb_entries_p0_d__T_1561_data; // @[tlb.scala 56:19]
  wire  _T_2377_v = _T_2376 ? tlb_entries_p1_v__T_1561_data : tlb_entries_p0_v__T_1561_data; // @[tlb.scala 56:19]
  wire  _T_2382 = ~_T_2377_v; // @[tlb.scala 59:18]
  wire  _T_2383 = ~_T_2377_d; // @[tlb.scala 63:25]
  wire  _T_2385 = _T_2383 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1507 = {{8'd0}, _T_2377_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2387 = _GEN_1507 & _T_1730; // @[tlb.scala 68:32]
  wire [43:0] _T_2388 = {_T_2387, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2393 = _T_2374 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2394 = _GEN_1461 & _T_2393; // @[tlb.scala 69:27]
  wire [43:0] _T_2395 = _T_2388 | _T_2394; // @[tlb.scala 70:29]
  wire [4:0] _GEN_292 = _T_2385 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_293 = _T_2385 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_294 = _T_2385 ? 44'h0 : _T_2395; // @[tlb.scala 63:53]
  wire [4:0] _GEN_295 = _T_2382 ? 5'h8 : _GEN_292; // @[tlb.scala 59:27]
  wire [4:0] _GEN_296 = _T_2382 ? _T_1989 : _GEN_293; // @[tlb.scala 59:27]
  wire [43:0] _GEN_297 = _T_2382 ? 44'h0 : _GEN_294; // @[tlb.scala 59:27]
  wire [31:0] _T_2399 = _T_1739 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2400 = {_T_2399, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2401 = _GEN_1461 & _T_2400; // @[tlb.scala 55:24]
  wire  _T_2402 = _T_2401 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2403_pfn = _T_2402 ? tlb_entries_p1_pfn__T_1562_data : tlb_entries_p0_pfn__T_1562_data; // @[tlb.scala 56:19]
  wire  _T_2403_d = _T_2402 ? tlb_entries_p1_d__T_1562_data : tlb_entries_p0_d__T_1562_data; // @[tlb.scala 56:19]
  wire  _T_2403_v = _T_2402 ? tlb_entries_p1_v__T_1562_data : tlb_entries_p0_v__T_1562_data; // @[tlb.scala 56:19]
  wire  _T_2408 = ~_T_2403_v; // @[tlb.scala 59:18]
  wire  _T_2409 = ~_T_2403_d; // @[tlb.scala 63:25]
  wire  _T_2411 = _T_2409 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1510 = {{8'd0}, _T_2403_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2413 = _GEN_1510 & _T_1740; // @[tlb.scala 68:32]
  wire [43:0] _T_2414 = {_T_2413, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2419 = _T_2400 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2420 = _GEN_1461 & _T_2419; // @[tlb.scala 69:27]
  wire [43:0] _T_2421 = _T_2414 | _T_2420; // @[tlb.scala 70:29]
  wire [4:0] _GEN_298 = _T_2411 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_299 = _T_2411 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_300 = _T_2411 ? 44'h0 : _T_2421; // @[tlb.scala 63:53]
  wire [4:0] _GEN_301 = _T_2408 ? 5'h8 : _GEN_298; // @[tlb.scala 59:27]
  wire [4:0] _GEN_302 = _T_2408 ? _T_1989 : _GEN_299; // @[tlb.scala 59:27]
  wire [43:0] _GEN_303 = _T_2408 ? 44'h0 : _GEN_300; // @[tlb.scala 59:27]
  wire [31:0] _T_2425 = _T_1749 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2426 = {_T_2425, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2427 = _GEN_1461 & _T_2426; // @[tlb.scala 55:24]
  wire  _T_2428 = _T_2427 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2429_pfn = _T_2428 ? tlb_entries_p1_pfn__T_1563_data : tlb_entries_p0_pfn__T_1563_data; // @[tlb.scala 56:19]
  wire  _T_2429_d = _T_2428 ? tlb_entries_p1_d__T_1563_data : tlb_entries_p0_d__T_1563_data; // @[tlb.scala 56:19]
  wire  _T_2429_v = _T_2428 ? tlb_entries_p1_v__T_1563_data : tlb_entries_p0_v__T_1563_data; // @[tlb.scala 56:19]
  wire  _T_2434 = ~_T_2429_v; // @[tlb.scala 59:18]
  wire  _T_2435 = ~_T_2429_d; // @[tlb.scala 63:25]
  wire  _T_2437 = _T_2435 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1513 = {{8'd0}, _T_2429_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2439 = _GEN_1513 & _T_1750; // @[tlb.scala 68:32]
  wire [43:0] _T_2440 = {_T_2439, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2445 = _T_2426 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2446 = _GEN_1461 & _T_2445; // @[tlb.scala 69:27]
  wire [43:0] _T_2447 = _T_2440 | _T_2446; // @[tlb.scala 70:29]
  wire [4:0] _GEN_304 = _T_2437 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_305 = _T_2437 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_306 = _T_2437 ? 44'h0 : _T_2447; // @[tlb.scala 63:53]
  wire [4:0] _GEN_307 = _T_2434 ? 5'h8 : _GEN_304; // @[tlb.scala 59:27]
  wire [4:0] _GEN_308 = _T_2434 ? _T_1989 : _GEN_305; // @[tlb.scala 59:27]
  wire [43:0] _GEN_309 = _T_2434 ? 44'h0 : _GEN_306; // @[tlb.scala 59:27]
  wire [31:0] _T_2451 = _T_1759 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2452 = {_T_2451, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2453 = _GEN_1461 & _T_2452; // @[tlb.scala 55:24]
  wire  _T_2454 = _T_2453 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2455_pfn = _T_2454 ? tlb_entries_p1_pfn__T_1564_data : tlb_entries_p0_pfn__T_1564_data; // @[tlb.scala 56:19]
  wire  _T_2455_d = _T_2454 ? tlb_entries_p1_d__T_1564_data : tlb_entries_p0_d__T_1564_data; // @[tlb.scala 56:19]
  wire  _T_2455_v = _T_2454 ? tlb_entries_p1_v__T_1564_data : tlb_entries_p0_v__T_1564_data; // @[tlb.scala 56:19]
  wire  _T_2460 = ~_T_2455_v; // @[tlb.scala 59:18]
  wire  _T_2461 = ~_T_2455_d; // @[tlb.scala 63:25]
  wire  _T_2463 = _T_2461 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1516 = {{8'd0}, _T_2455_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2465 = _GEN_1516 & _T_1760; // @[tlb.scala 68:32]
  wire [43:0] _T_2466 = {_T_2465, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2471 = _T_2452 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2472 = _GEN_1461 & _T_2471; // @[tlb.scala 69:27]
  wire [43:0] _T_2473 = _T_2466 | _T_2472; // @[tlb.scala 70:29]
  wire [4:0] _GEN_310 = _T_2463 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_311 = _T_2463 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_312 = _T_2463 ? 44'h0 : _T_2473; // @[tlb.scala 63:53]
  wire [4:0] _GEN_313 = _T_2460 ? 5'h8 : _GEN_310; // @[tlb.scala 59:27]
  wire [4:0] _GEN_314 = _T_2460 ? _T_1989 : _GEN_311; // @[tlb.scala 59:27]
  wire [43:0] _GEN_315 = _T_2460 ? 44'h0 : _GEN_312; // @[tlb.scala 59:27]
  wire [31:0] _T_2477 = _T_1769 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2478 = {_T_2477, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2479 = _GEN_1461 & _T_2478; // @[tlb.scala 55:24]
  wire  _T_2480 = _T_2479 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2481_pfn = _T_2480 ? tlb_entries_p1_pfn__T_1565_data : tlb_entries_p0_pfn__T_1565_data; // @[tlb.scala 56:19]
  wire  _T_2481_d = _T_2480 ? tlb_entries_p1_d__T_1565_data : tlb_entries_p0_d__T_1565_data; // @[tlb.scala 56:19]
  wire  _T_2481_v = _T_2480 ? tlb_entries_p1_v__T_1565_data : tlb_entries_p0_v__T_1565_data; // @[tlb.scala 56:19]
  wire  _T_2486 = ~_T_2481_v; // @[tlb.scala 59:18]
  wire  _T_2487 = ~_T_2481_d; // @[tlb.scala 63:25]
  wire  _T_2489 = _T_2487 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1519 = {{8'd0}, _T_2481_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2491 = _GEN_1519 & _T_1770; // @[tlb.scala 68:32]
  wire [43:0] _T_2492 = {_T_2491, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2497 = _T_2478 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2498 = _GEN_1461 & _T_2497; // @[tlb.scala 69:27]
  wire [43:0] _T_2499 = _T_2492 | _T_2498; // @[tlb.scala 70:29]
  wire [4:0] _GEN_316 = _T_2489 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_317 = _T_2489 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_318 = _T_2489 ? 44'h0 : _T_2499; // @[tlb.scala 63:53]
  wire [4:0] _GEN_319 = _T_2486 ? 5'h8 : _GEN_316; // @[tlb.scala 59:27]
  wire [4:0] _GEN_320 = _T_2486 ? _T_1989 : _GEN_317; // @[tlb.scala 59:27]
  wire [43:0] _GEN_321 = _T_2486 ? 44'h0 : _GEN_318; // @[tlb.scala 59:27]
  wire [31:0] _T_2503 = _T_1779 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2504 = {_T_2503, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2505 = _GEN_1461 & _T_2504; // @[tlb.scala 55:24]
  wire  _T_2506 = _T_2505 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2507_pfn = _T_2506 ? tlb_entries_p1_pfn__T_1566_data : tlb_entries_p0_pfn__T_1566_data; // @[tlb.scala 56:19]
  wire  _T_2507_d = _T_2506 ? tlb_entries_p1_d__T_1566_data : tlb_entries_p0_d__T_1566_data; // @[tlb.scala 56:19]
  wire  _T_2507_v = _T_2506 ? tlb_entries_p1_v__T_1566_data : tlb_entries_p0_v__T_1566_data; // @[tlb.scala 56:19]
  wire  _T_2512 = ~_T_2507_v; // @[tlb.scala 59:18]
  wire  _T_2513 = ~_T_2507_d; // @[tlb.scala 63:25]
  wire  _T_2515 = _T_2513 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1522 = {{8'd0}, _T_2507_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2517 = _GEN_1522 & _T_1780; // @[tlb.scala 68:32]
  wire [43:0] _T_2518 = {_T_2517, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2523 = _T_2504 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2524 = _GEN_1461 & _T_2523; // @[tlb.scala 69:27]
  wire [43:0] _T_2525 = _T_2518 | _T_2524; // @[tlb.scala 70:29]
  wire [4:0] _GEN_322 = _T_2515 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_323 = _T_2515 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_324 = _T_2515 ? 44'h0 : _T_2525; // @[tlb.scala 63:53]
  wire [4:0] _GEN_325 = _T_2512 ? 5'h8 : _GEN_322; // @[tlb.scala 59:27]
  wire [4:0] _GEN_326 = _T_2512 ? _T_1989 : _GEN_323; // @[tlb.scala 59:27]
  wire [43:0] _GEN_327 = _T_2512 ? 44'h0 : _GEN_324; // @[tlb.scala 59:27]
  wire [31:0] _T_2529 = _T_1789 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2530 = {_T_2529, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2531 = _GEN_1461 & _T_2530; // @[tlb.scala 55:24]
  wire  _T_2532 = _T_2531 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2533_pfn = _T_2532 ? tlb_entries_p1_pfn__T_1567_data : tlb_entries_p0_pfn__T_1567_data; // @[tlb.scala 56:19]
  wire  _T_2533_d = _T_2532 ? tlb_entries_p1_d__T_1567_data : tlb_entries_p0_d__T_1567_data; // @[tlb.scala 56:19]
  wire  _T_2533_v = _T_2532 ? tlb_entries_p1_v__T_1567_data : tlb_entries_p0_v__T_1567_data; // @[tlb.scala 56:19]
  wire  _T_2538 = ~_T_2533_v; // @[tlb.scala 59:18]
  wire  _T_2539 = ~_T_2533_d; // @[tlb.scala 63:25]
  wire  _T_2541 = _T_2539 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1525 = {{8'd0}, _T_2533_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2543 = _GEN_1525 & _T_1790; // @[tlb.scala 68:32]
  wire [43:0] _T_2544 = {_T_2543, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2549 = _T_2530 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2550 = _GEN_1461 & _T_2549; // @[tlb.scala 69:27]
  wire [43:0] _T_2551 = _T_2544 | _T_2550; // @[tlb.scala 70:29]
  wire [4:0] _GEN_328 = _T_2541 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_329 = _T_2541 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_330 = _T_2541 ? 44'h0 : _T_2551; // @[tlb.scala 63:53]
  wire [4:0] _GEN_331 = _T_2538 ? 5'h8 : _GEN_328; // @[tlb.scala 59:27]
  wire [4:0] _GEN_332 = _T_2538 ? _T_1989 : _GEN_329; // @[tlb.scala 59:27]
  wire [43:0] _GEN_333 = _T_2538 ? 44'h0 : _GEN_330; // @[tlb.scala 59:27]
  wire [31:0] _T_2555 = _T_1799 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2556 = {_T_2555, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2557 = _GEN_1461 & _T_2556; // @[tlb.scala 55:24]
  wire  _T_2558 = _T_2557 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2559_pfn = _T_2558 ? tlb_entries_p1_pfn__T_1568_data : tlb_entries_p0_pfn__T_1568_data; // @[tlb.scala 56:19]
  wire  _T_2559_d = _T_2558 ? tlb_entries_p1_d__T_1568_data : tlb_entries_p0_d__T_1568_data; // @[tlb.scala 56:19]
  wire  _T_2559_v = _T_2558 ? tlb_entries_p1_v__T_1568_data : tlb_entries_p0_v__T_1568_data; // @[tlb.scala 56:19]
  wire  _T_2564 = ~_T_2559_v; // @[tlb.scala 59:18]
  wire  _T_2565 = ~_T_2559_d; // @[tlb.scala 63:25]
  wire  _T_2567 = _T_2565 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1528 = {{8'd0}, _T_2559_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2569 = _GEN_1528 & _T_1800; // @[tlb.scala 68:32]
  wire [43:0] _T_2570 = {_T_2569, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2575 = _T_2556 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2576 = _GEN_1461 & _T_2575; // @[tlb.scala 69:27]
  wire [43:0] _T_2577 = _T_2570 | _T_2576; // @[tlb.scala 70:29]
  wire [4:0] _GEN_334 = _T_2567 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_335 = _T_2567 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_336 = _T_2567 ? 44'h0 : _T_2577; // @[tlb.scala 63:53]
  wire [4:0] _GEN_337 = _T_2564 ? 5'h8 : _GEN_334; // @[tlb.scala 59:27]
  wire [4:0] _GEN_338 = _T_2564 ? _T_1989 : _GEN_335; // @[tlb.scala 59:27]
  wire [43:0] _GEN_339 = _T_2564 ? 44'h0 : _GEN_336; // @[tlb.scala 59:27]
  wire [31:0] _T_2581 = _T_1809 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2582 = {_T_2581, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2583 = _GEN_1461 & _T_2582; // @[tlb.scala 55:24]
  wire  _T_2584 = _T_2583 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2585_pfn = _T_2584 ? tlb_entries_p1_pfn__T_1569_data : tlb_entries_p0_pfn__T_1569_data; // @[tlb.scala 56:19]
  wire  _T_2585_d = _T_2584 ? tlb_entries_p1_d__T_1569_data : tlb_entries_p0_d__T_1569_data; // @[tlb.scala 56:19]
  wire  _T_2585_v = _T_2584 ? tlb_entries_p1_v__T_1569_data : tlb_entries_p0_v__T_1569_data; // @[tlb.scala 56:19]
  wire  _T_2590 = ~_T_2585_v; // @[tlb.scala 59:18]
  wire  _T_2591 = ~_T_2585_d; // @[tlb.scala 63:25]
  wire  _T_2593 = _T_2591 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1531 = {{8'd0}, _T_2585_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2595 = _GEN_1531 & _T_1810; // @[tlb.scala 68:32]
  wire [43:0] _T_2596 = {_T_2595, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2601 = _T_2582 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2602 = _GEN_1461 & _T_2601; // @[tlb.scala 69:27]
  wire [43:0] _T_2603 = _T_2596 | _T_2602; // @[tlb.scala 70:29]
  wire [4:0] _GEN_340 = _T_2593 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_341 = _T_2593 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_342 = _T_2593 ? 44'h0 : _T_2603; // @[tlb.scala 63:53]
  wire [4:0] _GEN_343 = _T_2590 ? 5'h8 : _GEN_340; // @[tlb.scala 59:27]
  wire [4:0] _GEN_344 = _T_2590 ? _T_1989 : _GEN_341; // @[tlb.scala 59:27]
  wire [43:0] _GEN_345 = _T_2590 ? 44'h0 : _GEN_342; // @[tlb.scala 59:27]
  wire [31:0] _T_2607 = _T_1819 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2608 = {_T_2607, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2609 = _GEN_1461 & _T_2608; // @[tlb.scala 55:24]
  wire  _T_2610 = _T_2609 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2611_pfn = _T_2610 ? tlb_entries_p1_pfn__T_1570_data : tlb_entries_p0_pfn__T_1570_data; // @[tlb.scala 56:19]
  wire  _T_2611_d = _T_2610 ? tlb_entries_p1_d__T_1570_data : tlb_entries_p0_d__T_1570_data; // @[tlb.scala 56:19]
  wire  _T_2611_v = _T_2610 ? tlb_entries_p1_v__T_1570_data : tlb_entries_p0_v__T_1570_data; // @[tlb.scala 56:19]
  wire  _T_2616 = ~_T_2611_v; // @[tlb.scala 59:18]
  wire  _T_2617 = ~_T_2611_d; // @[tlb.scala 63:25]
  wire  _T_2619 = _T_2617 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1534 = {{8'd0}, _T_2611_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2621 = _GEN_1534 & _T_1820; // @[tlb.scala 68:32]
  wire [43:0] _T_2622 = {_T_2621, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2627 = _T_2608 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2628 = _GEN_1461 & _T_2627; // @[tlb.scala 69:27]
  wire [43:0] _T_2629 = _T_2622 | _T_2628; // @[tlb.scala 70:29]
  wire [4:0] _GEN_346 = _T_2619 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_347 = _T_2619 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_348 = _T_2619 ? 44'h0 : _T_2629; // @[tlb.scala 63:53]
  wire [4:0] _GEN_349 = _T_2616 ? 5'h8 : _GEN_346; // @[tlb.scala 59:27]
  wire [4:0] _GEN_350 = _T_2616 ? _T_1989 : _GEN_347; // @[tlb.scala 59:27]
  wire [43:0] _GEN_351 = _T_2616 ? 44'h0 : _GEN_348; // @[tlb.scala 59:27]
  wire [31:0] _T_2633 = _T_1829 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2634 = {_T_2633, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2635 = _GEN_1461 & _T_2634; // @[tlb.scala 55:24]
  wire  _T_2636 = _T_2635 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2637_pfn = _T_2636 ? tlb_entries_p1_pfn__T_1571_data : tlb_entries_p0_pfn__T_1571_data; // @[tlb.scala 56:19]
  wire  _T_2637_d = _T_2636 ? tlb_entries_p1_d__T_1571_data : tlb_entries_p0_d__T_1571_data; // @[tlb.scala 56:19]
  wire  _T_2637_v = _T_2636 ? tlb_entries_p1_v__T_1571_data : tlb_entries_p0_v__T_1571_data; // @[tlb.scala 56:19]
  wire  _T_2642 = ~_T_2637_v; // @[tlb.scala 59:18]
  wire  _T_2643 = ~_T_2637_d; // @[tlb.scala 63:25]
  wire  _T_2645 = _T_2643 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1537 = {{8'd0}, _T_2637_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2647 = _GEN_1537 & _T_1830; // @[tlb.scala 68:32]
  wire [43:0] _T_2648 = {_T_2647, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2653 = _T_2634 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2654 = _GEN_1461 & _T_2653; // @[tlb.scala 69:27]
  wire [43:0] _T_2655 = _T_2648 | _T_2654; // @[tlb.scala 70:29]
  wire [4:0] _GEN_352 = _T_2645 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_353 = _T_2645 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_354 = _T_2645 ? 44'h0 : _T_2655; // @[tlb.scala 63:53]
  wire [4:0] _GEN_355 = _T_2642 ? 5'h8 : _GEN_352; // @[tlb.scala 59:27]
  wire [4:0] _GEN_356 = _T_2642 ? _T_1989 : _GEN_353; // @[tlb.scala 59:27]
  wire [43:0] _GEN_357 = _T_2642 ? 44'h0 : _GEN_354; // @[tlb.scala 59:27]
  wire [31:0] _T_2659 = _T_1839 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2660 = {_T_2659, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2661 = _GEN_1461 & _T_2660; // @[tlb.scala 55:24]
  wire  _T_2662 = _T_2661 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2663_pfn = _T_2662 ? tlb_entries_p1_pfn__T_1572_data : tlb_entries_p0_pfn__T_1572_data; // @[tlb.scala 56:19]
  wire  _T_2663_d = _T_2662 ? tlb_entries_p1_d__T_1572_data : tlb_entries_p0_d__T_1572_data; // @[tlb.scala 56:19]
  wire  _T_2663_v = _T_2662 ? tlb_entries_p1_v__T_1572_data : tlb_entries_p0_v__T_1572_data; // @[tlb.scala 56:19]
  wire  _T_2668 = ~_T_2663_v; // @[tlb.scala 59:18]
  wire  _T_2669 = ~_T_2663_d; // @[tlb.scala 63:25]
  wire  _T_2671 = _T_2669 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1540 = {{8'd0}, _T_2663_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2673 = _GEN_1540 & _T_1840; // @[tlb.scala 68:32]
  wire [43:0] _T_2674 = {_T_2673, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2679 = _T_2660 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2680 = _GEN_1461 & _T_2679; // @[tlb.scala 69:27]
  wire [43:0] _T_2681 = _T_2674 | _T_2680; // @[tlb.scala 70:29]
  wire [4:0] _GEN_358 = _T_2671 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_359 = _T_2671 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_360 = _T_2671 ? 44'h0 : _T_2681; // @[tlb.scala 63:53]
  wire [4:0] _GEN_361 = _T_2668 ? 5'h8 : _GEN_358; // @[tlb.scala 59:27]
  wire [4:0] _GEN_362 = _T_2668 ? _T_1989 : _GEN_359; // @[tlb.scala 59:27]
  wire [43:0] _GEN_363 = _T_2668 ? 44'h0 : _GEN_360; // @[tlb.scala 59:27]
  wire [31:0] _T_2685 = _T_1849 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2686 = {_T_2685, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2687 = _GEN_1461 & _T_2686; // @[tlb.scala 55:24]
  wire  _T_2688 = _T_2687 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2689_pfn = _T_2688 ? tlb_entries_p1_pfn__T_1573_data : tlb_entries_p0_pfn__T_1573_data; // @[tlb.scala 56:19]
  wire  _T_2689_d = _T_2688 ? tlb_entries_p1_d__T_1573_data : tlb_entries_p0_d__T_1573_data; // @[tlb.scala 56:19]
  wire  _T_2689_v = _T_2688 ? tlb_entries_p1_v__T_1573_data : tlb_entries_p0_v__T_1573_data; // @[tlb.scala 56:19]
  wire  _T_2694 = ~_T_2689_v; // @[tlb.scala 59:18]
  wire  _T_2695 = ~_T_2689_d; // @[tlb.scala 63:25]
  wire  _T_2697 = _T_2695 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1543 = {{8'd0}, _T_2689_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2699 = _GEN_1543 & _T_1850; // @[tlb.scala 68:32]
  wire [43:0] _T_2700 = {_T_2699, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2705 = _T_2686 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2706 = _GEN_1461 & _T_2705; // @[tlb.scala 69:27]
  wire [43:0] _T_2707 = _T_2700 | _T_2706; // @[tlb.scala 70:29]
  wire [4:0] _GEN_364 = _T_2697 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_365 = _T_2697 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_366 = _T_2697 ? 44'h0 : _T_2707; // @[tlb.scala 63:53]
  wire [4:0] _GEN_367 = _T_2694 ? 5'h8 : _GEN_364; // @[tlb.scala 59:27]
  wire [4:0] _GEN_368 = _T_2694 ? _T_1989 : _GEN_365; // @[tlb.scala 59:27]
  wire [43:0] _GEN_369 = _T_2694 ? 44'h0 : _GEN_366; // @[tlb.scala 59:27]
  wire [31:0] _T_2711 = _T_1859 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2712 = {_T_2711, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2713 = _GEN_1461 & _T_2712; // @[tlb.scala 55:24]
  wire  _T_2714 = _T_2713 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2715_pfn = _T_2714 ? tlb_entries_p1_pfn__T_1574_data : tlb_entries_p0_pfn__T_1574_data; // @[tlb.scala 56:19]
  wire  _T_2715_d = _T_2714 ? tlb_entries_p1_d__T_1574_data : tlb_entries_p0_d__T_1574_data; // @[tlb.scala 56:19]
  wire  _T_2715_v = _T_2714 ? tlb_entries_p1_v__T_1574_data : tlb_entries_p0_v__T_1574_data; // @[tlb.scala 56:19]
  wire  _T_2720 = ~_T_2715_v; // @[tlb.scala 59:18]
  wire  _T_2721 = ~_T_2715_d; // @[tlb.scala 63:25]
  wire  _T_2723 = _T_2721 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1546 = {{8'd0}, _T_2715_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2725 = _GEN_1546 & _T_1860; // @[tlb.scala 68:32]
  wire [43:0] _T_2726 = {_T_2725, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2731 = _T_2712 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2732 = _GEN_1461 & _T_2731; // @[tlb.scala 69:27]
  wire [43:0] _T_2733 = _T_2726 | _T_2732; // @[tlb.scala 70:29]
  wire [4:0] _GEN_370 = _T_2723 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_371 = _T_2723 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_372 = _T_2723 ? 44'h0 : _T_2733; // @[tlb.scala 63:53]
  wire [4:0] _GEN_373 = _T_2720 ? 5'h8 : _GEN_370; // @[tlb.scala 59:27]
  wire [4:0] _GEN_374 = _T_2720 ? _T_1989 : _GEN_371; // @[tlb.scala 59:27]
  wire [43:0] _GEN_375 = _T_2720 ? 44'h0 : _GEN_372; // @[tlb.scala 59:27]
  wire [31:0] _T_2737 = _T_1869 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2738 = {_T_2737, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2739 = _GEN_1461 & _T_2738; // @[tlb.scala 55:24]
  wire  _T_2740 = _T_2739 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2741_pfn = _T_2740 ? tlb_entries_p1_pfn__T_1575_data : tlb_entries_p0_pfn__T_1575_data; // @[tlb.scala 56:19]
  wire  _T_2741_d = _T_2740 ? tlb_entries_p1_d__T_1575_data : tlb_entries_p0_d__T_1575_data; // @[tlb.scala 56:19]
  wire  _T_2741_v = _T_2740 ? tlb_entries_p1_v__T_1575_data : tlb_entries_p0_v__T_1575_data; // @[tlb.scala 56:19]
  wire  _T_2746 = ~_T_2741_v; // @[tlb.scala 59:18]
  wire  _T_2747 = ~_T_2741_d; // @[tlb.scala 63:25]
  wire  _T_2749 = _T_2747 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1549 = {{8'd0}, _T_2741_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2751 = _GEN_1549 & _T_1870; // @[tlb.scala 68:32]
  wire [43:0] _T_2752 = {_T_2751, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2757 = _T_2738 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2758 = _GEN_1461 & _T_2757; // @[tlb.scala 69:27]
  wire [43:0] _T_2759 = _T_2752 | _T_2758; // @[tlb.scala 70:29]
  wire [4:0] _GEN_376 = _T_2749 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_377 = _T_2749 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_378 = _T_2749 ? 44'h0 : _T_2759; // @[tlb.scala 63:53]
  wire [4:0] _GEN_379 = _T_2746 ? 5'h8 : _GEN_376; // @[tlb.scala 59:27]
  wire [4:0] _GEN_380 = _T_2746 ? _T_1989 : _GEN_377; // @[tlb.scala 59:27]
  wire [43:0] _GEN_381 = _T_2746 ? 44'h0 : _GEN_378; // @[tlb.scala 59:27]
  wire [31:0] _T_2763 = _T_1879 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2764 = {_T_2763, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2765 = _GEN_1461 & _T_2764; // @[tlb.scala 55:24]
  wire  _T_2766 = _T_2765 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2767_pfn = _T_2766 ? tlb_entries_p1_pfn__T_1576_data : tlb_entries_p0_pfn__T_1576_data; // @[tlb.scala 56:19]
  wire  _T_2767_d = _T_2766 ? tlb_entries_p1_d__T_1576_data : tlb_entries_p0_d__T_1576_data; // @[tlb.scala 56:19]
  wire  _T_2767_v = _T_2766 ? tlb_entries_p1_v__T_1576_data : tlb_entries_p0_v__T_1576_data; // @[tlb.scala 56:19]
  wire  _T_2772 = ~_T_2767_v; // @[tlb.scala 59:18]
  wire  _T_2773 = ~_T_2767_d; // @[tlb.scala 63:25]
  wire  _T_2775 = _T_2773 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1552 = {{8'd0}, _T_2767_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2777 = _GEN_1552 & _T_1880; // @[tlb.scala 68:32]
  wire [43:0] _T_2778 = {_T_2777, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2783 = _T_2764 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2784 = _GEN_1461 & _T_2783; // @[tlb.scala 69:27]
  wire [43:0] _T_2785 = _T_2778 | _T_2784; // @[tlb.scala 70:29]
  wire [4:0] _GEN_382 = _T_2775 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_383 = _T_2775 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_384 = _T_2775 ? 44'h0 : _T_2785; // @[tlb.scala 63:53]
  wire [4:0] _GEN_385 = _T_2772 ? 5'h8 : _GEN_382; // @[tlb.scala 59:27]
  wire [4:0] _GEN_386 = _T_2772 ? _T_1989 : _GEN_383; // @[tlb.scala 59:27]
  wire [43:0] _GEN_387 = _T_2772 ? 44'h0 : _GEN_384; // @[tlb.scala 59:27]
  wire [31:0] _T_2789 = _T_1889 + 32'h1; // @[tlb.scala 55:33]
  wire [43:0] _T_2790 = {_T_2789, 12'h0}; // @[tlb.scala 55:40]
  wire [43:0] _T_2791 = _GEN_1461 & _T_2790; // @[tlb.scala 55:24]
  wire  _T_2792 = _T_2791 != 44'h0; // @[tlb.scala 55:48]
  wire [23:0] _T_2793_pfn = _T_2792 ? tlb_entries_p1_pfn__T_1577_data : tlb_entries_p0_pfn__T_1577_data; // @[tlb.scala 56:19]
  wire  _T_2793_d = _T_2792 ? tlb_entries_p1_d__T_1577_data : tlb_entries_p0_d__T_1577_data; // @[tlb.scala 56:19]
  wire  _T_2793_v = _T_2792 ? tlb_entries_p1_v__T_1577_data : tlb_entries_p0_v__T_1577_data; // @[tlb.scala 56:19]
  wire  _T_2798 = ~_T_2793_v; // @[tlb.scala 59:18]
  wire  _T_2799 = ~_T_2793_d; // @[tlb.scala 63:25]
  wire  _T_2801 = _T_2799 & _T_1544_func; // @[tlb.scala 63:33]
  wire [31:0] _GEN_1555 = {{8'd0}, _T_2793_pfn}; // @[tlb.scala 68:32]
  wire [31:0] _T_2803 = _GEN_1555 & _T_1890; // @[tlb.scala 68:32]
  wire [43:0] _T_2804 = {_T_2803, 12'h0}; // @[tlb.scala 68:41]
  wire [43:0] _T_2809 = _T_2790 - 44'h1; // @[tlb.scala 69:51]
  wire [43:0] _T_2810 = _GEN_1461 & _T_2809; // @[tlb.scala 69:27]
  wire [43:0] _T_2811 = _T_2804 | _T_2810; // @[tlb.scala 70:29]
  wire [4:0] _GEN_388 = _T_2801 ? 5'h9 : 5'h0; // @[tlb.scala 63:53]
  wire [4:0] _GEN_389 = _T_2801 ? 5'h1 : _T_1989; // @[tlb.scala 63:53]
  wire [43:0] _GEN_390 = _T_2801 ? 44'h0 : _T_2811; // @[tlb.scala 63:53]
  wire [4:0] _GEN_391 = _T_2798 ? 5'h8 : _GEN_388; // @[tlb.scala 59:27]
  wire [4:0] _GEN_392 = _T_2798 ? _T_1989 : _GEN_389; // @[tlb.scala 59:27]
  wire [43:0] _GEN_393 = _T_2798 ? 44'h0 : _GEN_390; // @[tlb.scala 59:27]
  wire [7:0] _T_1991_ex_asid = tlb_entries_asid__T_1546_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2815 = {_GEN_205,_GEN_206,_T_1544_vaddr,_T_1991_ex_asid,_GEN_207[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2816 = _T_1977[0] ? _T_2815 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2017_ex_asid = tlb_entries_asid__T_1547_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2820 = {_GEN_211,_GEN_212,_T_1544_vaddr,_T_2017_ex_asid,_GEN_213[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2821 = _T_1977[1] ? _T_2820 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2043_ex_asid = tlb_entries_asid__T_1548_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2825 = {_GEN_217,_GEN_218,_T_1544_vaddr,_T_2043_ex_asid,_GEN_219[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2826 = _T_1977[2] ? _T_2825 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2069_ex_asid = tlb_entries_asid__T_1549_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2830 = {_GEN_223,_GEN_224,_T_1544_vaddr,_T_2069_ex_asid,_GEN_225[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2831 = _T_1977[3] ? _T_2830 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2095_ex_asid = tlb_entries_asid__T_1550_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2835 = {_GEN_229,_GEN_230,_T_1544_vaddr,_T_2095_ex_asid,_GEN_231[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2836 = _T_1977[4] ? _T_2835 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2121_ex_asid = tlb_entries_asid__T_1551_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2840 = {_GEN_235,_GEN_236,_T_1544_vaddr,_T_2121_ex_asid,_GEN_237[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2841 = _T_1977[5] ? _T_2840 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2147_ex_asid = tlb_entries_asid__T_1552_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2845 = {_GEN_241,_GEN_242,_T_1544_vaddr,_T_2147_ex_asid,_GEN_243[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2846 = _T_1977[6] ? _T_2845 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2173_ex_asid = tlb_entries_asid__T_1553_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2850 = {_GEN_247,_GEN_248,_T_1544_vaddr,_T_2173_ex_asid,_GEN_249[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2851 = _T_1977[7] ? _T_2850 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2199_ex_asid = tlb_entries_asid__T_1554_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2855 = {_GEN_253,_GEN_254,_T_1544_vaddr,_T_2199_ex_asid,_GEN_255[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2856 = _T_1977[8] ? _T_2855 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2225_ex_asid = tlb_entries_asid__T_1555_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2860 = {_GEN_259,_GEN_260,_T_1544_vaddr,_T_2225_ex_asid,_GEN_261[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2861 = _T_1977[9] ? _T_2860 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2251_ex_asid = tlb_entries_asid__T_1556_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2865 = {_GEN_265,_GEN_266,_T_1544_vaddr,_T_2251_ex_asid,_GEN_267[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2866 = _T_1977[10] ? _T_2865 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2277_ex_asid = tlb_entries_asid__T_1557_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2870 = {_GEN_271,_GEN_272,_T_1544_vaddr,_T_2277_ex_asid,_GEN_273[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2871 = _T_1977[11] ? _T_2870 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2303_ex_asid = tlb_entries_asid__T_1558_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2875 = {_GEN_277,_GEN_278,_T_1544_vaddr,_T_2303_ex_asid,_GEN_279[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2876 = _T_1977[12] ? _T_2875 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2329_ex_asid = tlb_entries_asid__T_1559_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2880 = {_GEN_283,_GEN_284,_T_1544_vaddr,_T_2329_ex_asid,_GEN_285[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2881 = _T_1977[13] ? _T_2880 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2355_ex_asid = tlb_entries_asid__T_1560_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2885 = {_GEN_289,_GEN_290,_T_1544_vaddr,_T_2355_ex_asid,_GEN_291[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2886 = _T_1977[14] ? _T_2885 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2381_ex_asid = tlb_entries_asid__T_1561_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2890 = {_GEN_295,_GEN_296,_T_1544_vaddr,_T_2381_ex_asid,_GEN_297[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2891 = _T_1977[15] ? _T_2890 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2407_ex_asid = tlb_entries_asid__T_1562_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2895 = {_GEN_301,_GEN_302,_T_1544_vaddr,_T_2407_ex_asid,_GEN_303[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2896 = _T_1977[16] ? _T_2895 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2433_ex_asid = tlb_entries_asid__T_1563_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2900 = {_GEN_307,_GEN_308,_T_1544_vaddr,_T_2433_ex_asid,_GEN_309[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2901 = _T_1977[17] ? _T_2900 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2459_ex_asid = tlb_entries_asid__T_1564_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2905 = {_GEN_313,_GEN_314,_T_1544_vaddr,_T_2459_ex_asid,_GEN_315[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2906 = _T_1977[18] ? _T_2905 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2485_ex_asid = tlb_entries_asid__T_1565_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2910 = {_GEN_319,_GEN_320,_T_1544_vaddr,_T_2485_ex_asid,_GEN_321[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2911 = _T_1977[19] ? _T_2910 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2511_ex_asid = tlb_entries_asid__T_1566_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2915 = {_GEN_325,_GEN_326,_T_1544_vaddr,_T_2511_ex_asid,_GEN_327[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2916 = _T_1977[20] ? _T_2915 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2537_ex_asid = tlb_entries_asid__T_1567_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2920 = {_GEN_331,_GEN_332,_T_1544_vaddr,_T_2537_ex_asid,_GEN_333[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2921 = _T_1977[21] ? _T_2920 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2563_ex_asid = tlb_entries_asid__T_1568_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2925 = {_GEN_337,_GEN_338,_T_1544_vaddr,_T_2563_ex_asid,_GEN_339[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2926 = _T_1977[22] ? _T_2925 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2589_ex_asid = tlb_entries_asid__T_1569_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2930 = {_GEN_343,_GEN_344,_T_1544_vaddr,_T_2589_ex_asid,_GEN_345[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2931 = _T_1977[23] ? _T_2930 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2615_ex_asid = tlb_entries_asid__T_1570_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2935 = {_GEN_349,_GEN_350,_T_1544_vaddr,_T_2615_ex_asid,_GEN_351[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2936 = _T_1977[24] ? _T_2935 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2641_ex_asid = tlb_entries_asid__T_1571_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2940 = {_GEN_355,_GEN_356,_T_1544_vaddr,_T_2641_ex_asid,_GEN_357[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2941 = _T_1977[25] ? _T_2940 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2667_ex_asid = tlb_entries_asid__T_1572_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2945 = {_GEN_361,_GEN_362,_T_1544_vaddr,_T_2667_ex_asid,_GEN_363[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2946 = _T_1977[26] ? _T_2945 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2693_ex_asid = tlb_entries_asid__T_1573_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2950 = {_GEN_367,_GEN_368,_T_1544_vaddr,_T_2693_ex_asid,_GEN_369[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2951 = _T_1977[27] ? _T_2950 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2719_ex_asid = tlb_entries_asid__T_1574_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2955 = {_GEN_373,_GEN_374,_T_1544_vaddr,_T_2719_ex_asid,_GEN_375[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2956 = _T_1977[28] ? _T_2955 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2745_ex_asid = tlb_entries_asid__T_1575_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2960 = {_GEN_379,_GEN_380,_T_1544_vaddr,_T_2745_ex_asid,_GEN_381[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2961 = _T_1977[29] ? _T_2960 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2771_ex_asid = tlb_entries_asid__T_1576_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2965 = {_GEN_385,_GEN_386,_T_1544_vaddr,_T_2771_ex_asid,_GEN_387[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2966 = _T_1977[30] ? _T_2965 : 82'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_2797_ex_asid = tlb_entries_asid__T_1577_data; // @[tlb.scala 74:17]
  wire [81:0] _T_2970 = {_GEN_391,_GEN_392,_T_1544_vaddr,_T_2797_ex_asid,_GEN_393[31:0]}; // @[Mux.scala 27:72]
  wire [81:0] _T_2971 = _T_1977[31] ? _T_2970 : 82'h0; // @[Mux.scala 27:72]
  wire [81:0] _T_2972 = _T_2816 | _T_2821; // @[Mux.scala 27:72]
  wire [81:0] _T_2973 = _T_2972 | _T_2826; // @[Mux.scala 27:72]
  wire [81:0] _T_2974 = _T_2973 | _T_2831; // @[Mux.scala 27:72]
  wire [81:0] _T_2975 = _T_2974 | _T_2836; // @[Mux.scala 27:72]
  wire [81:0] _T_2976 = _T_2975 | _T_2841; // @[Mux.scala 27:72]
  wire [81:0] _T_2977 = _T_2976 | _T_2846; // @[Mux.scala 27:72]
  wire [81:0] _T_2978 = _T_2977 | _T_2851; // @[Mux.scala 27:72]
  wire [81:0] _T_2979 = _T_2978 | _T_2856; // @[Mux.scala 27:72]
  wire [81:0] _T_2980 = _T_2979 | _T_2861; // @[Mux.scala 27:72]
  wire [81:0] _T_2981 = _T_2980 | _T_2866; // @[Mux.scala 27:72]
  wire [81:0] _T_2982 = _T_2981 | _T_2871; // @[Mux.scala 27:72]
  wire [81:0] _T_2983 = _T_2982 | _T_2876; // @[Mux.scala 27:72]
  wire [81:0] _T_2984 = _T_2983 | _T_2881; // @[Mux.scala 27:72]
  wire [81:0] _T_2985 = _T_2984 | _T_2886; // @[Mux.scala 27:72]
  wire [81:0] _T_2986 = _T_2985 | _T_2891; // @[Mux.scala 27:72]
  wire [81:0] _T_2987 = _T_2986 | _T_2896; // @[Mux.scala 27:72]
  wire [81:0] _T_2988 = _T_2987 | _T_2901; // @[Mux.scala 27:72]
  wire [81:0] _T_2989 = _T_2988 | _T_2906; // @[Mux.scala 27:72]
  wire [81:0] _T_2990 = _T_2989 | _T_2911; // @[Mux.scala 27:72]
  wire [81:0] _T_2991 = _T_2990 | _T_2916; // @[Mux.scala 27:72]
  wire [81:0] _T_2992 = _T_2991 | _T_2921; // @[Mux.scala 27:72]
  wire [81:0] _T_2993 = _T_2992 | _T_2926; // @[Mux.scala 27:72]
  wire [81:0] _T_2994 = _T_2993 | _T_2931; // @[Mux.scala 27:72]
  wire [81:0] _T_2995 = _T_2994 | _T_2936; // @[Mux.scala 27:72]
  wire [81:0] _T_2996 = _T_2995 | _T_2941; // @[Mux.scala 27:72]
  wire [81:0] _T_2997 = _T_2996 | _T_2946; // @[Mux.scala 27:72]
  wire [81:0] _T_2998 = _T_2997 | _T_2951; // @[Mux.scala 27:72]
  wire [81:0] _T_2999 = _T_2998 | _T_2956; // @[Mux.scala 27:72]
  wire [81:0] _T_3000 = _T_2999 | _T_2961; // @[Mux.scala 27:72]
  wire [81:0] _T_3001 = _T_3000 | _T_2966; // @[Mux.scala 27:72]
  wire [81:0] _T_3002 = _T_3001 | _T_2971; // @[Mux.scala 27:72]
  wire [4:0] _T_3014_ex_et = _T_1979 ? 5'h7 : _T_3002[81:77]; // @[tlb.scala 102:8]
  wire [4:0] _T_3014_ex_code = _T_1979 ? _T_1989 : _T_3002[76:72]; // @[tlb.scala 102:8]
  wire [7:0] _T_3014_ex_asid = _T_1979 ? 8'h0 : _T_3002[39:32]; // @[tlb.scala 102:8]
  wire [31:0] _T_3014_paddr = _T_1979 ? 32'h0 : _T_3002[31:0]; // @[tlb.scala 102:8]
  wire  _T_3016 = _T_1544_vaddr[31:29] == 3'h4; // @[tlb.scala 111:12]
  wire  _T_3017 = _T_1544_vaddr[31:29] == 3'h5; // @[tlb.scala 111:27]
  wire  _T_3018 = _T_3016 | _T_3017; // @[tlb.scala 111:20]
  wire [29:0] _T_3020 = {1'h0,_T_1544_vaddr[28:0]}; // @[Cat.scala 29:58]
  wire  _T_3021 = _T_1544_vaddr[31:29] == 3'h6; // @[tlb.scala 112:12]
  wire [29:0] _T_3023 = {1'h0,_T_3014_paddr[28:0]}; // @[Cat.scala 29:58]
  wire  _T_3024 = _T_1544_vaddr[31:29] == 3'h7; // @[tlb.scala 113:12]
  wire  _T_3026 = ~_T_1544_vaddr[31]; // @[tlb.scala 114:15]
  wire [31:0] _T_3029 = io_status_ERL ? _T_1544_vaddr : {{2'd0}, _T_3023}; // @[tlb.scala 114:30]
  wire [29:0] _T_3030 = _T_3018 ? _T_3020 : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_3031 = _T_3021 ? _T_3023 : 30'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_3032 = _T_3024 ? _T_1544_vaddr : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_3033 = _T_3026 ? _T_3029 : 32'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_3034 = _T_3030 | _T_3031; // @[Mux.scala 27:72]
  wire [31:0] _GEN_1557 = {{2'd0}, _T_3034}; // @[Mux.scala 27:72]
  wire [31:0] _T_3035 = _GEN_1557 | _T_3032; // @[Mux.scala 27:72]
  wire [4:0] _T_3044 = io_status_ERL ? 5'h0 : _T_3014_ex_et; // @[tlb.scala 120:30]
  wire [4:0] _T_3046 = _T_3021 ? _T_3014_ex_et : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3047 = _T_3026 ? _T_3044 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3049 = _T_3046 | _T_3047; // @[Mux.scala 27:72]
  wire [1:0] _T_3054 = _T_1544_is_aligned ? _T_1544_vaddr[1:0] : 2'h0; // @[tlb.scala 148:23]
  wire  _T_3056 = _T_1544_len == 2'h1; // @[tlb.scala 152:22]
  wire  _T_3058 = _T_1544_len == 2'h3; // @[tlb.scala 153:22]
  wire  _T_3059 = _T_3054 != 2'h0; // @[tlb.scala 153:45]
  wire  _T_3061 = _T_3056 & _T_3054[0]; // @[Mux.scala 27:72]
  wire  _T_3062 = _T_3058 & _T_3059; // @[Mux.scala 27:72]
  wire  _T_3064 = _T_3061 | _T_3062; // @[Mux.scala 27:72]
  wire [4:0] _T_3069 = _T_1988 ? 5'h4 : 5'h5; // @[tlb.scala 157:24]
  wire  _T_3080 = ~io_ex_flush_valid; // @[tlb.scala 168:18]
  wire  _T_3083 = 5'h0 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3084 = 5'h1 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3085 = 5'h2 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3086 = 5'h3 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3087 = 5'h4 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3088 = 5'h5 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3089 = 5'h6 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3090 = 5'h7 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3091 = 5'h8 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3092 = 5'h9 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3093 = 5'ha == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3094 = 5'hb == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3095 = 5'hc == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3096 = 5'hd == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3097 = 5'he == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3098 = 5'hf == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3099 = 5'h10 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3100 = 5'h11 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3101 = 5'h12 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3102 = 5'h13 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3103 = 5'h14 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3104 = 5'h15 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3105 = 5'h16 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3106 = 5'h17 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3107 = 5'h18 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3108 = 5'h19 == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3109 = 5'h1a == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3110 = 5'h1b == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3111 = 5'h1c == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3112 = 5'h1d == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3113 = 5'h1e == io_rport_index; // @[tlb.scala 192:10]
  wire  _T_3114 = 5'h1f == io_rport_index; // @[tlb.scala 192:10]
  wire [30:0] _T_3119 = {tlb_entries_p0_d_tlb_entry_ports_0_r_data,tlb_entries_p0_v_tlb_entry_ports_0_r_data,tlb_entries_p1_pfn_tlb_entry_ports_0_r_data,tlb_entries_p1_c_tlb_entry_ports_0_r_data,tlb_entries_p1_d_tlb_entry_ports_0_r_data,tlb_entries_p1_v_tlb_entry_ports_0_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3125 = {tlb_entries_pagemask_tlb_entry_ports_0_r_data,tlb_entries_vpn_tlb_entry_ports_0_r_data,tlb_entries_g_tlb_entry_ports_0_r_data,tlb_entries_asid_tlb_entry_ports_0_r_data,tlb_entries_p0_pfn_tlb_entry_ports_0_r_data,tlb_entries_p0_c_tlb_entry_ports_0_r_data,_T_3119}; // @[Mux.scala 27:72]
  wire [101:0] _T_3126 = _T_3083 ? _T_3125 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3131 = {tlb_entries_p0_d_tlb_entry_ports_1_r_data,tlb_entries_p0_v_tlb_entry_ports_1_r_data,tlb_entries_p1_pfn_tlb_entry_ports_1_r_data,tlb_entries_p1_c_tlb_entry_ports_1_r_data,tlb_entries_p1_d_tlb_entry_ports_1_r_data,tlb_entries_p1_v_tlb_entry_ports_1_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3137 = {tlb_entries_pagemask_tlb_entry_ports_1_r_data,tlb_entries_vpn_tlb_entry_ports_1_r_data,tlb_entries_g_tlb_entry_ports_1_r_data,tlb_entries_asid_tlb_entry_ports_1_r_data,tlb_entries_p0_pfn_tlb_entry_ports_1_r_data,tlb_entries_p0_c_tlb_entry_ports_1_r_data,_T_3131}; // @[Mux.scala 27:72]
  wire [101:0] _T_3138 = _T_3084 ? _T_3137 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3143 = {tlb_entries_p0_d_tlb_entry_ports_2_r_data,tlb_entries_p0_v_tlb_entry_ports_2_r_data,tlb_entries_p1_pfn_tlb_entry_ports_2_r_data,tlb_entries_p1_c_tlb_entry_ports_2_r_data,tlb_entries_p1_d_tlb_entry_ports_2_r_data,tlb_entries_p1_v_tlb_entry_ports_2_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3149 = {tlb_entries_pagemask_tlb_entry_ports_2_r_data,tlb_entries_vpn_tlb_entry_ports_2_r_data,tlb_entries_g_tlb_entry_ports_2_r_data,tlb_entries_asid_tlb_entry_ports_2_r_data,tlb_entries_p0_pfn_tlb_entry_ports_2_r_data,tlb_entries_p0_c_tlb_entry_ports_2_r_data,_T_3143}; // @[Mux.scala 27:72]
  wire [101:0] _T_3150 = _T_3085 ? _T_3149 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3155 = {tlb_entries_p0_d_tlb_entry_ports_3_r_data,tlb_entries_p0_v_tlb_entry_ports_3_r_data,tlb_entries_p1_pfn_tlb_entry_ports_3_r_data,tlb_entries_p1_c_tlb_entry_ports_3_r_data,tlb_entries_p1_d_tlb_entry_ports_3_r_data,tlb_entries_p1_v_tlb_entry_ports_3_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3161 = {tlb_entries_pagemask_tlb_entry_ports_3_r_data,tlb_entries_vpn_tlb_entry_ports_3_r_data,tlb_entries_g_tlb_entry_ports_3_r_data,tlb_entries_asid_tlb_entry_ports_3_r_data,tlb_entries_p0_pfn_tlb_entry_ports_3_r_data,tlb_entries_p0_c_tlb_entry_ports_3_r_data,_T_3155}; // @[Mux.scala 27:72]
  wire [101:0] _T_3162 = _T_3086 ? _T_3161 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3167 = {tlb_entries_p0_d_tlb_entry_ports_4_r_data,tlb_entries_p0_v_tlb_entry_ports_4_r_data,tlb_entries_p1_pfn_tlb_entry_ports_4_r_data,tlb_entries_p1_c_tlb_entry_ports_4_r_data,tlb_entries_p1_d_tlb_entry_ports_4_r_data,tlb_entries_p1_v_tlb_entry_ports_4_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3173 = {tlb_entries_pagemask_tlb_entry_ports_4_r_data,tlb_entries_vpn_tlb_entry_ports_4_r_data,tlb_entries_g_tlb_entry_ports_4_r_data,tlb_entries_asid_tlb_entry_ports_4_r_data,tlb_entries_p0_pfn_tlb_entry_ports_4_r_data,tlb_entries_p0_c_tlb_entry_ports_4_r_data,_T_3167}; // @[Mux.scala 27:72]
  wire [101:0] _T_3174 = _T_3087 ? _T_3173 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3179 = {tlb_entries_p0_d_tlb_entry_ports_5_r_data,tlb_entries_p0_v_tlb_entry_ports_5_r_data,tlb_entries_p1_pfn_tlb_entry_ports_5_r_data,tlb_entries_p1_c_tlb_entry_ports_5_r_data,tlb_entries_p1_d_tlb_entry_ports_5_r_data,tlb_entries_p1_v_tlb_entry_ports_5_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3185 = {tlb_entries_pagemask_tlb_entry_ports_5_r_data,tlb_entries_vpn_tlb_entry_ports_5_r_data,tlb_entries_g_tlb_entry_ports_5_r_data,tlb_entries_asid_tlb_entry_ports_5_r_data,tlb_entries_p0_pfn_tlb_entry_ports_5_r_data,tlb_entries_p0_c_tlb_entry_ports_5_r_data,_T_3179}; // @[Mux.scala 27:72]
  wire [101:0] _T_3186 = _T_3088 ? _T_3185 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3191 = {tlb_entries_p0_d_tlb_entry_ports_6_r_data,tlb_entries_p0_v_tlb_entry_ports_6_r_data,tlb_entries_p1_pfn_tlb_entry_ports_6_r_data,tlb_entries_p1_c_tlb_entry_ports_6_r_data,tlb_entries_p1_d_tlb_entry_ports_6_r_data,tlb_entries_p1_v_tlb_entry_ports_6_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3197 = {tlb_entries_pagemask_tlb_entry_ports_6_r_data,tlb_entries_vpn_tlb_entry_ports_6_r_data,tlb_entries_g_tlb_entry_ports_6_r_data,tlb_entries_asid_tlb_entry_ports_6_r_data,tlb_entries_p0_pfn_tlb_entry_ports_6_r_data,tlb_entries_p0_c_tlb_entry_ports_6_r_data,_T_3191}; // @[Mux.scala 27:72]
  wire [101:0] _T_3198 = _T_3089 ? _T_3197 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3203 = {tlb_entries_p0_d_tlb_entry_ports_7_r_data,tlb_entries_p0_v_tlb_entry_ports_7_r_data,tlb_entries_p1_pfn_tlb_entry_ports_7_r_data,tlb_entries_p1_c_tlb_entry_ports_7_r_data,tlb_entries_p1_d_tlb_entry_ports_7_r_data,tlb_entries_p1_v_tlb_entry_ports_7_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3209 = {tlb_entries_pagemask_tlb_entry_ports_7_r_data,tlb_entries_vpn_tlb_entry_ports_7_r_data,tlb_entries_g_tlb_entry_ports_7_r_data,tlb_entries_asid_tlb_entry_ports_7_r_data,tlb_entries_p0_pfn_tlb_entry_ports_7_r_data,tlb_entries_p0_c_tlb_entry_ports_7_r_data,_T_3203}; // @[Mux.scala 27:72]
  wire [101:0] _T_3210 = _T_3090 ? _T_3209 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3215 = {tlb_entries_p0_d_tlb_entry_ports_8_r_data,tlb_entries_p0_v_tlb_entry_ports_8_r_data,tlb_entries_p1_pfn_tlb_entry_ports_8_r_data,tlb_entries_p1_c_tlb_entry_ports_8_r_data,tlb_entries_p1_d_tlb_entry_ports_8_r_data,tlb_entries_p1_v_tlb_entry_ports_8_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3221 = {tlb_entries_pagemask_tlb_entry_ports_8_r_data,tlb_entries_vpn_tlb_entry_ports_8_r_data,tlb_entries_g_tlb_entry_ports_8_r_data,tlb_entries_asid_tlb_entry_ports_8_r_data,tlb_entries_p0_pfn_tlb_entry_ports_8_r_data,tlb_entries_p0_c_tlb_entry_ports_8_r_data,_T_3215}; // @[Mux.scala 27:72]
  wire [101:0] _T_3222 = _T_3091 ? _T_3221 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3227 = {tlb_entries_p0_d_tlb_entry_ports_9_r_data,tlb_entries_p0_v_tlb_entry_ports_9_r_data,tlb_entries_p1_pfn_tlb_entry_ports_9_r_data,tlb_entries_p1_c_tlb_entry_ports_9_r_data,tlb_entries_p1_d_tlb_entry_ports_9_r_data,tlb_entries_p1_v_tlb_entry_ports_9_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3233 = {tlb_entries_pagemask_tlb_entry_ports_9_r_data,tlb_entries_vpn_tlb_entry_ports_9_r_data,tlb_entries_g_tlb_entry_ports_9_r_data,tlb_entries_asid_tlb_entry_ports_9_r_data,tlb_entries_p0_pfn_tlb_entry_ports_9_r_data,tlb_entries_p0_c_tlb_entry_ports_9_r_data,_T_3227}; // @[Mux.scala 27:72]
  wire [101:0] _T_3234 = _T_3092 ? _T_3233 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3239 = {tlb_entries_p0_d_tlb_entry_ports_10_r_data,tlb_entries_p0_v_tlb_entry_ports_10_r_data,tlb_entries_p1_pfn_tlb_entry_ports_10_r_data,tlb_entries_p1_c_tlb_entry_ports_10_r_data,tlb_entries_p1_d_tlb_entry_ports_10_r_data,tlb_entries_p1_v_tlb_entry_ports_10_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3245 = {tlb_entries_pagemask_tlb_entry_ports_10_r_data,tlb_entries_vpn_tlb_entry_ports_10_r_data,tlb_entries_g_tlb_entry_ports_10_r_data,tlb_entries_asid_tlb_entry_ports_10_r_data,tlb_entries_p0_pfn_tlb_entry_ports_10_r_data,tlb_entries_p0_c_tlb_entry_ports_10_r_data,_T_3239}; // @[Mux.scala 27:72]
  wire [101:0] _T_3246 = _T_3093 ? _T_3245 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3251 = {tlb_entries_p0_d_tlb_entry_ports_11_r_data,tlb_entries_p0_v_tlb_entry_ports_11_r_data,tlb_entries_p1_pfn_tlb_entry_ports_11_r_data,tlb_entries_p1_c_tlb_entry_ports_11_r_data,tlb_entries_p1_d_tlb_entry_ports_11_r_data,tlb_entries_p1_v_tlb_entry_ports_11_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3257 = {tlb_entries_pagemask_tlb_entry_ports_11_r_data,tlb_entries_vpn_tlb_entry_ports_11_r_data,tlb_entries_g_tlb_entry_ports_11_r_data,tlb_entries_asid_tlb_entry_ports_11_r_data,tlb_entries_p0_pfn_tlb_entry_ports_11_r_data,tlb_entries_p0_c_tlb_entry_ports_11_r_data,_T_3251}; // @[Mux.scala 27:72]
  wire [101:0] _T_3258 = _T_3094 ? _T_3257 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3263 = {tlb_entries_p0_d_tlb_entry_ports_12_r_data,tlb_entries_p0_v_tlb_entry_ports_12_r_data,tlb_entries_p1_pfn_tlb_entry_ports_12_r_data,tlb_entries_p1_c_tlb_entry_ports_12_r_data,tlb_entries_p1_d_tlb_entry_ports_12_r_data,tlb_entries_p1_v_tlb_entry_ports_12_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3269 = {tlb_entries_pagemask_tlb_entry_ports_12_r_data,tlb_entries_vpn_tlb_entry_ports_12_r_data,tlb_entries_g_tlb_entry_ports_12_r_data,tlb_entries_asid_tlb_entry_ports_12_r_data,tlb_entries_p0_pfn_tlb_entry_ports_12_r_data,tlb_entries_p0_c_tlb_entry_ports_12_r_data,_T_3263}; // @[Mux.scala 27:72]
  wire [101:0] _T_3270 = _T_3095 ? _T_3269 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3275 = {tlb_entries_p0_d_tlb_entry_ports_13_r_data,tlb_entries_p0_v_tlb_entry_ports_13_r_data,tlb_entries_p1_pfn_tlb_entry_ports_13_r_data,tlb_entries_p1_c_tlb_entry_ports_13_r_data,tlb_entries_p1_d_tlb_entry_ports_13_r_data,tlb_entries_p1_v_tlb_entry_ports_13_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3281 = {tlb_entries_pagemask_tlb_entry_ports_13_r_data,tlb_entries_vpn_tlb_entry_ports_13_r_data,tlb_entries_g_tlb_entry_ports_13_r_data,tlb_entries_asid_tlb_entry_ports_13_r_data,tlb_entries_p0_pfn_tlb_entry_ports_13_r_data,tlb_entries_p0_c_tlb_entry_ports_13_r_data,_T_3275}; // @[Mux.scala 27:72]
  wire [101:0] _T_3282 = _T_3096 ? _T_3281 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3287 = {tlb_entries_p0_d_tlb_entry_ports_14_r_data,tlb_entries_p0_v_tlb_entry_ports_14_r_data,tlb_entries_p1_pfn_tlb_entry_ports_14_r_data,tlb_entries_p1_c_tlb_entry_ports_14_r_data,tlb_entries_p1_d_tlb_entry_ports_14_r_data,tlb_entries_p1_v_tlb_entry_ports_14_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3293 = {tlb_entries_pagemask_tlb_entry_ports_14_r_data,tlb_entries_vpn_tlb_entry_ports_14_r_data,tlb_entries_g_tlb_entry_ports_14_r_data,tlb_entries_asid_tlb_entry_ports_14_r_data,tlb_entries_p0_pfn_tlb_entry_ports_14_r_data,tlb_entries_p0_c_tlb_entry_ports_14_r_data,_T_3287}; // @[Mux.scala 27:72]
  wire [101:0] _T_3294 = _T_3097 ? _T_3293 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3299 = {tlb_entries_p0_d_tlb_entry_ports_15_r_data,tlb_entries_p0_v_tlb_entry_ports_15_r_data,tlb_entries_p1_pfn_tlb_entry_ports_15_r_data,tlb_entries_p1_c_tlb_entry_ports_15_r_data,tlb_entries_p1_d_tlb_entry_ports_15_r_data,tlb_entries_p1_v_tlb_entry_ports_15_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3305 = {tlb_entries_pagemask_tlb_entry_ports_15_r_data,tlb_entries_vpn_tlb_entry_ports_15_r_data,tlb_entries_g_tlb_entry_ports_15_r_data,tlb_entries_asid_tlb_entry_ports_15_r_data,tlb_entries_p0_pfn_tlb_entry_ports_15_r_data,tlb_entries_p0_c_tlb_entry_ports_15_r_data,_T_3299}; // @[Mux.scala 27:72]
  wire [101:0] _T_3306 = _T_3098 ? _T_3305 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3311 = {tlb_entries_p0_d_tlb_entry_ports_16_r_data,tlb_entries_p0_v_tlb_entry_ports_16_r_data,tlb_entries_p1_pfn_tlb_entry_ports_16_r_data,tlb_entries_p1_c_tlb_entry_ports_16_r_data,tlb_entries_p1_d_tlb_entry_ports_16_r_data,tlb_entries_p1_v_tlb_entry_ports_16_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3317 = {tlb_entries_pagemask_tlb_entry_ports_16_r_data,tlb_entries_vpn_tlb_entry_ports_16_r_data,tlb_entries_g_tlb_entry_ports_16_r_data,tlb_entries_asid_tlb_entry_ports_16_r_data,tlb_entries_p0_pfn_tlb_entry_ports_16_r_data,tlb_entries_p0_c_tlb_entry_ports_16_r_data,_T_3311}; // @[Mux.scala 27:72]
  wire [101:0] _T_3318 = _T_3099 ? _T_3317 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3323 = {tlb_entries_p0_d_tlb_entry_ports_17_r_data,tlb_entries_p0_v_tlb_entry_ports_17_r_data,tlb_entries_p1_pfn_tlb_entry_ports_17_r_data,tlb_entries_p1_c_tlb_entry_ports_17_r_data,tlb_entries_p1_d_tlb_entry_ports_17_r_data,tlb_entries_p1_v_tlb_entry_ports_17_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3329 = {tlb_entries_pagemask_tlb_entry_ports_17_r_data,tlb_entries_vpn_tlb_entry_ports_17_r_data,tlb_entries_g_tlb_entry_ports_17_r_data,tlb_entries_asid_tlb_entry_ports_17_r_data,tlb_entries_p0_pfn_tlb_entry_ports_17_r_data,tlb_entries_p0_c_tlb_entry_ports_17_r_data,_T_3323}; // @[Mux.scala 27:72]
  wire [101:0] _T_3330 = _T_3100 ? _T_3329 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3335 = {tlb_entries_p0_d_tlb_entry_ports_18_r_data,tlb_entries_p0_v_tlb_entry_ports_18_r_data,tlb_entries_p1_pfn_tlb_entry_ports_18_r_data,tlb_entries_p1_c_tlb_entry_ports_18_r_data,tlb_entries_p1_d_tlb_entry_ports_18_r_data,tlb_entries_p1_v_tlb_entry_ports_18_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3341 = {tlb_entries_pagemask_tlb_entry_ports_18_r_data,tlb_entries_vpn_tlb_entry_ports_18_r_data,tlb_entries_g_tlb_entry_ports_18_r_data,tlb_entries_asid_tlb_entry_ports_18_r_data,tlb_entries_p0_pfn_tlb_entry_ports_18_r_data,tlb_entries_p0_c_tlb_entry_ports_18_r_data,_T_3335}; // @[Mux.scala 27:72]
  wire [101:0] _T_3342 = _T_3101 ? _T_3341 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3347 = {tlb_entries_p0_d_tlb_entry_ports_19_r_data,tlb_entries_p0_v_tlb_entry_ports_19_r_data,tlb_entries_p1_pfn_tlb_entry_ports_19_r_data,tlb_entries_p1_c_tlb_entry_ports_19_r_data,tlb_entries_p1_d_tlb_entry_ports_19_r_data,tlb_entries_p1_v_tlb_entry_ports_19_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3353 = {tlb_entries_pagemask_tlb_entry_ports_19_r_data,tlb_entries_vpn_tlb_entry_ports_19_r_data,tlb_entries_g_tlb_entry_ports_19_r_data,tlb_entries_asid_tlb_entry_ports_19_r_data,tlb_entries_p0_pfn_tlb_entry_ports_19_r_data,tlb_entries_p0_c_tlb_entry_ports_19_r_data,_T_3347}; // @[Mux.scala 27:72]
  wire [101:0] _T_3354 = _T_3102 ? _T_3353 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3359 = {tlb_entries_p0_d_tlb_entry_ports_20_r_data,tlb_entries_p0_v_tlb_entry_ports_20_r_data,tlb_entries_p1_pfn_tlb_entry_ports_20_r_data,tlb_entries_p1_c_tlb_entry_ports_20_r_data,tlb_entries_p1_d_tlb_entry_ports_20_r_data,tlb_entries_p1_v_tlb_entry_ports_20_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3365 = {tlb_entries_pagemask_tlb_entry_ports_20_r_data,tlb_entries_vpn_tlb_entry_ports_20_r_data,tlb_entries_g_tlb_entry_ports_20_r_data,tlb_entries_asid_tlb_entry_ports_20_r_data,tlb_entries_p0_pfn_tlb_entry_ports_20_r_data,tlb_entries_p0_c_tlb_entry_ports_20_r_data,_T_3359}; // @[Mux.scala 27:72]
  wire [101:0] _T_3366 = _T_3103 ? _T_3365 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3371 = {tlb_entries_p0_d_tlb_entry_ports_21_r_data,tlb_entries_p0_v_tlb_entry_ports_21_r_data,tlb_entries_p1_pfn_tlb_entry_ports_21_r_data,tlb_entries_p1_c_tlb_entry_ports_21_r_data,tlb_entries_p1_d_tlb_entry_ports_21_r_data,tlb_entries_p1_v_tlb_entry_ports_21_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3377 = {tlb_entries_pagemask_tlb_entry_ports_21_r_data,tlb_entries_vpn_tlb_entry_ports_21_r_data,tlb_entries_g_tlb_entry_ports_21_r_data,tlb_entries_asid_tlb_entry_ports_21_r_data,tlb_entries_p0_pfn_tlb_entry_ports_21_r_data,tlb_entries_p0_c_tlb_entry_ports_21_r_data,_T_3371}; // @[Mux.scala 27:72]
  wire [101:0] _T_3378 = _T_3104 ? _T_3377 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3383 = {tlb_entries_p0_d_tlb_entry_ports_22_r_data,tlb_entries_p0_v_tlb_entry_ports_22_r_data,tlb_entries_p1_pfn_tlb_entry_ports_22_r_data,tlb_entries_p1_c_tlb_entry_ports_22_r_data,tlb_entries_p1_d_tlb_entry_ports_22_r_data,tlb_entries_p1_v_tlb_entry_ports_22_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3389 = {tlb_entries_pagemask_tlb_entry_ports_22_r_data,tlb_entries_vpn_tlb_entry_ports_22_r_data,tlb_entries_g_tlb_entry_ports_22_r_data,tlb_entries_asid_tlb_entry_ports_22_r_data,tlb_entries_p0_pfn_tlb_entry_ports_22_r_data,tlb_entries_p0_c_tlb_entry_ports_22_r_data,_T_3383}; // @[Mux.scala 27:72]
  wire [101:0] _T_3390 = _T_3105 ? _T_3389 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3395 = {tlb_entries_p0_d_tlb_entry_ports_23_r_data,tlb_entries_p0_v_tlb_entry_ports_23_r_data,tlb_entries_p1_pfn_tlb_entry_ports_23_r_data,tlb_entries_p1_c_tlb_entry_ports_23_r_data,tlb_entries_p1_d_tlb_entry_ports_23_r_data,tlb_entries_p1_v_tlb_entry_ports_23_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3401 = {tlb_entries_pagemask_tlb_entry_ports_23_r_data,tlb_entries_vpn_tlb_entry_ports_23_r_data,tlb_entries_g_tlb_entry_ports_23_r_data,tlb_entries_asid_tlb_entry_ports_23_r_data,tlb_entries_p0_pfn_tlb_entry_ports_23_r_data,tlb_entries_p0_c_tlb_entry_ports_23_r_data,_T_3395}; // @[Mux.scala 27:72]
  wire [101:0] _T_3402 = _T_3106 ? _T_3401 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3407 = {tlb_entries_p0_d_tlb_entry_ports_24_r_data,tlb_entries_p0_v_tlb_entry_ports_24_r_data,tlb_entries_p1_pfn_tlb_entry_ports_24_r_data,tlb_entries_p1_c_tlb_entry_ports_24_r_data,tlb_entries_p1_d_tlb_entry_ports_24_r_data,tlb_entries_p1_v_tlb_entry_ports_24_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3413 = {tlb_entries_pagemask_tlb_entry_ports_24_r_data,tlb_entries_vpn_tlb_entry_ports_24_r_data,tlb_entries_g_tlb_entry_ports_24_r_data,tlb_entries_asid_tlb_entry_ports_24_r_data,tlb_entries_p0_pfn_tlb_entry_ports_24_r_data,tlb_entries_p0_c_tlb_entry_ports_24_r_data,_T_3407}; // @[Mux.scala 27:72]
  wire [101:0] _T_3414 = _T_3107 ? _T_3413 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3419 = {tlb_entries_p0_d_tlb_entry_ports_25_r_data,tlb_entries_p0_v_tlb_entry_ports_25_r_data,tlb_entries_p1_pfn_tlb_entry_ports_25_r_data,tlb_entries_p1_c_tlb_entry_ports_25_r_data,tlb_entries_p1_d_tlb_entry_ports_25_r_data,tlb_entries_p1_v_tlb_entry_ports_25_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3425 = {tlb_entries_pagemask_tlb_entry_ports_25_r_data,tlb_entries_vpn_tlb_entry_ports_25_r_data,tlb_entries_g_tlb_entry_ports_25_r_data,tlb_entries_asid_tlb_entry_ports_25_r_data,tlb_entries_p0_pfn_tlb_entry_ports_25_r_data,tlb_entries_p0_c_tlb_entry_ports_25_r_data,_T_3419}; // @[Mux.scala 27:72]
  wire [101:0] _T_3426 = _T_3108 ? _T_3425 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3431 = {tlb_entries_p0_d_tlb_entry_ports_26_r_data,tlb_entries_p0_v_tlb_entry_ports_26_r_data,tlb_entries_p1_pfn_tlb_entry_ports_26_r_data,tlb_entries_p1_c_tlb_entry_ports_26_r_data,tlb_entries_p1_d_tlb_entry_ports_26_r_data,tlb_entries_p1_v_tlb_entry_ports_26_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3437 = {tlb_entries_pagemask_tlb_entry_ports_26_r_data,tlb_entries_vpn_tlb_entry_ports_26_r_data,tlb_entries_g_tlb_entry_ports_26_r_data,tlb_entries_asid_tlb_entry_ports_26_r_data,tlb_entries_p0_pfn_tlb_entry_ports_26_r_data,tlb_entries_p0_c_tlb_entry_ports_26_r_data,_T_3431}; // @[Mux.scala 27:72]
  wire [101:0] _T_3438 = _T_3109 ? _T_3437 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3443 = {tlb_entries_p0_d_tlb_entry_ports_27_r_data,tlb_entries_p0_v_tlb_entry_ports_27_r_data,tlb_entries_p1_pfn_tlb_entry_ports_27_r_data,tlb_entries_p1_c_tlb_entry_ports_27_r_data,tlb_entries_p1_d_tlb_entry_ports_27_r_data,tlb_entries_p1_v_tlb_entry_ports_27_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3449 = {tlb_entries_pagemask_tlb_entry_ports_27_r_data,tlb_entries_vpn_tlb_entry_ports_27_r_data,tlb_entries_g_tlb_entry_ports_27_r_data,tlb_entries_asid_tlb_entry_ports_27_r_data,tlb_entries_p0_pfn_tlb_entry_ports_27_r_data,tlb_entries_p0_c_tlb_entry_ports_27_r_data,_T_3443}; // @[Mux.scala 27:72]
  wire [101:0] _T_3450 = _T_3110 ? _T_3449 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3455 = {tlb_entries_p0_d_tlb_entry_ports_28_r_data,tlb_entries_p0_v_tlb_entry_ports_28_r_data,tlb_entries_p1_pfn_tlb_entry_ports_28_r_data,tlb_entries_p1_c_tlb_entry_ports_28_r_data,tlb_entries_p1_d_tlb_entry_ports_28_r_data,tlb_entries_p1_v_tlb_entry_ports_28_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3461 = {tlb_entries_pagemask_tlb_entry_ports_28_r_data,tlb_entries_vpn_tlb_entry_ports_28_r_data,tlb_entries_g_tlb_entry_ports_28_r_data,tlb_entries_asid_tlb_entry_ports_28_r_data,tlb_entries_p0_pfn_tlb_entry_ports_28_r_data,tlb_entries_p0_c_tlb_entry_ports_28_r_data,_T_3455}; // @[Mux.scala 27:72]
  wire [101:0] _T_3462 = _T_3111 ? _T_3461 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3467 = {tlb_entries_p0_d_tlb_entry_ports_29_r_data,tlb_entries_p0_v_tlb_entry_ports_29_r_data,tlb_entries_p1_pfn_tlb_entry_ports_29_r_data,tlb_entries_p1_c_tlb_entry_ports_29_r_data,tlb_entries_p1_d_tlb_entry_ports_29_r_data,tlb_entries_p1_v_tlb_entry_ports_29_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3473 = {tlb_entries_pagemask_tlb_entry_ports_29_r_data,tlb_entries_vpn_tlb_entry_ports_29_r_data,tlb_entries_g_tlb_entry_ports_29_r_data,tlb_entries_asid_tlb_entry_ports_29_r_data,tlb_entries_p0_pfn_tlb_entry_ports_29_r_data,tlb_entries_p0_c_tlb_entry_ports_29_r_data,_T_3467}; // @[Mux.scala 27:72]
  wire [101:0] _T_3474 = _T_3112 ? _T_3473 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3479 = {tlb_entries_p0_d_tlb_entry_ports_30_r_data,tlb_entries_p0_v_tlb_entry_ports_30_r_data,tlb_entries_p1_pfn_tlb_entry_ports_30_r_data,tlb_entries_p1_c_tlb_entry_ports_30_r_data,tlb_entries_p1_d_tlb_entry_ports_30_r_data,tlb_entries_p1_v_tlb_entry_ports_30_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3485 = {tlb_entries_pagemask_tlb_entry_ports_30_r_data,tlb_entries_vpn_tlb_entry_ports_30_r_data,tlb_entries_g_tlb_entry_ports_30_r_data,tlb_entries_asid_tlb_entry_ports_30_r_data,tlb_entries_p0_pfn_tlb_entry_ports_30_r_data,tlb_entries_p0_c_tlb_entry_ports_30_r_data,_T_3479}; // @[Mux.scala 27:72]
  wire [101:0] _T_3486 = _T_3113 ? _T_3485 : 102'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_3491 = {tlb_entries_p0_d_tlb_entry_ports_31_r_data,tlb_entries_p0_v_tlb_entry_ports_31_r_data,tlb_entries_p1_pfn_tlb_entry_ports_31_r_data,tlb_entries_p1_c_tlb_entry_ports_31_r_data,tlb_entries_p1_d_tlb_entry_ports_31_r_data,tlb_entries_p1_v_tlb_entry_ports_31_r_data}; // @[Mux.scala 27:72]
  wire [101:0] _T_3497 = {tlb_entries_pagemask_tlb_entry_ports_31_r_data,tlb_entries_vpn_tlb_entry_ports_31_r_data,tlb_entries_g_tlb_entry_ports_31_r_data,tlb_entries_asid_tlb_entry_ports_31_r_data,tlb_entries_p0_pfn_tlb_entry_ports_31_r_data,tlb_entries_p0_c_tlb_entry_ports_31_r_data,_T_3491}; // @[Mux.scala 27:72]
  wire [101:0] _T_3498 = _T_3114 ? _T_3497 : 102'h0; // @[Mux.scala 27:72]
  wire [101:0] _T_3499 = _T_3126 | _T_3138; // @[Mux.scala 27:72]
  wire [101:0] _T_3500 = _T_3499 | _T_3150; // @[Mux.scala 27:72]
  wire [101:0] _T_3501 = _T_3500 | _T_3162; // @[Mux.scala 27:72]
  wire [101:0] _T_3502 = _T_3501 | _T_3174; // @[Mux.scala 27:72]
  wire [101:0] _T_3503 = _T_3502 | _T_3186; // @[Mux.scala 27:72]
  wire [101:0] _T_3504 = _T_3503 | _T_3198; // @[Mux.scala 27:72]
  wire [101:0] _T_3505 = _T_3504 | _T_3210; // @[Mux.scala 27:72]
  wire [101:0] _T_3506 = _T_3505 | _T_3222; // @[Mux.scala 27:72]
  wire [101:0] _T_3507 = _T_3506 | _T_3234; // @[Mux.scala 27:72]
  wire [101:0] _T_3508 = _T_3507 | _T_3246; // @[Mux.scala 27:72]
  wire [101:0] _T_3509 = _T_3508 | _T_3258; // @[Mux.scala 27:72]
  wire [101:0] _T_3510 = _T_3509 | _T_3270; // @[Mux.scala 27:72]
  wire [101:0] _T_3511 = _T_3510 | _T_3282; // @[Mux.scala 27:72]
  wire [101:0] _T_3512 = _T_3511 | _T_3294; // @[Mux.scala 27:72]
  wire [101:0] _T_3513 = _T_3512 | _T_3306; // @[Mux.scala 27:72]
  wire [101:0] _T_3514 = _T_3513 | _T_3318; // @[Mux.scala 27:72]
  wire [101:0] _T_3515 = _T_3514 | _T_3330; // @[Mux.scala 27:72]
  wire [101:0] _T_3516 = _T_3515 | _T_3342; // @[Mux.scala 27:72]
  wire [101:0] _T_3517 = _T_3516 | _T_3354; // @[Mux.scala 27:72]
  wire [101:0] _T_3518 = _T_3517 | _T_3366; // @[Mux.scala 27:72]
  wire [101:0] _T_3519 = _T_3518 | _T_3378; // @[Mux.scala 27:72]
  wire [101:0] _T_3520 = _T_3519 | _T_3390; // @[Mux.scala 27:72]
  wire [101:0] _T_3521 = _T_3520 | _T_3402; // @[Mux.scala 27:72]
  wire [101:0] _T_3522 = _T_3521 | _T_3414; // @[Mux.scala 27:72]
  wire [101:0] _T_3523 = _T_3522 | _T_3426; // @[Mux.scala 27:72]
  wire [101:0] _T_3524 = _T_3523 | _T_3438; // @[Mux.scala 27:72]
  wire [101:0] _T_3525 = _T_3524 | _T_3450; // @[Mux.scala 27:72]
  wire [101:0] _T_3526 = _T_3525 | _T_3462; // @[Mux.scala 27:72]
  wire [101:0] _T_3527 = _T_3526 | _T_3474; // @[Mux.scala 27:72]
  wire [101:0] _T_3528 = _T_3527 | _T_3486; // @[Mux.scala 27:72]
  wire [101:0] _T_3529 = _T_3528 | _T_3498; // @[Mux.scala 27:72]
  wire  _T_3545 = io_wport_valid & _T_3080; // @[tlb.scala 193:24]
  wire  _T_3546 = 5'h0 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3547 = 5'h1 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3548 = 5'h2 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3549 = 5'h3 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3550 = 5'h4 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3551 = 5'h5 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3552 = 5'h6 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3553 = 5'h7 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3554 = 5'h8 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3555 = 5'h9 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3556 = 5'ha == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3557 = 5'hb == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3558 = 5'hc == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3559 = 5'hd == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3560 = 5'he == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3561 = 5'hf == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3562 = 5'h10 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3563 = 5'h11 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3564 = 5'h12 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3565 = 5'h13 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3566 = 5'h14 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3567 = 5'h15 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3568 = 5'h16 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3569 = 5'h17 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3570 = 5'h18 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3571 = 5'h19 == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3572 = 5'h1a == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3573 = 5'h1b == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3574 = 5'h1c == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3575 = 5'h1d == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3576 = 5'h1e == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _T_3577 = 5'h1f == io_wport_bits_index; // @[tlb.scala 195:17]
  wire  _GEN_813 = _T_3545 & _T_3546; // @[tlb.scala 193:47]
  wire  _GEN_826 = _T_3545 & _T_3547; // @[tlb.scala 193:47]
  wire  _GEN_839 = _T_3545 & _T_3548; // @[tlb.scala 193:47]
  wire  _GEN_852 = _T_3545 & _T_3549; // @[tlb.scala 193:47]
  wire  _GEN_865 = _T_3545 & _T_3550; // @[tlb.scala 193:47]
  wire  _GEN_878 = _T_3545 & _T_3551; // @[tlb.scala 193:47]
  wire  _GEN_891 = _T_3545 & _T_3552; // @[tlb.scala 193:47]
  wire  _GEN_904 = _T_3545 & _T_3553; // @[tlb.scala 193:47]
  wire  _GEN_917 = _T_3545 & _T_3554; // @[tlb.scala 193:47]
  wire  _GEN_930 = _T_3545 & _T_3555; // @[tlb.scala 193:47]
  wire  _GEN_943 = _T_3545 & _T_3556; // @[tlb.scala 193:47]
  wire  _GEN_956 = _T_3545 & _T_3557; // @[tlb.scala 193:47]
  wire  _GEN_969 = _T_3545 & _T_3558; // @[tlb.scala 193:47]
  wire  _GEN_982 = _T_3545 & _T_3559; // @[tlb.scala 193:47]
  wire  _GEN_995 = _T_3545 & _T_3560; // @[tlb.scala 193:47]
  wire  _GEN_1008 = _T_3545 & _T_3561; // @[tlb.scala 193:47]
  wire  _GEN_1021 = _T_3545 & _T_3562; // @[tlb.scala 193:47]
  wire  _GEN_1034 = _T_3545 & _T_3563; // @[tlb.scala 193:47]
  wire  _GEN_1047 = _T_3545 & _T_3564; // @[tlb.scala 193:47]
  wire  _GEN_1060 = _T_3545 & _T_3565; // @[tlb.scala 193:47]
  wire  _GEN_1073 = _T_3545 & _T_3566; // @[tlb.scala 193:47]
  wire  _GEN_1086 = _T_3545 & _T_3567; // @[tlb.scala 193:47]
  wire  _GEN_1099 = _T_3545 & _T_3568; // @[tlb.scala 193:47]
  wire  _GEN_1112 = _T_3545 & _T_3569; // @[tlb.scala 193:47]
  wire  _GEN_1125 = _T_3545 & _T_3570; // @[tlb.scala 193:47]
  wire  _GEN_1138 = _T_3545 & _T_3571; // @[tlb.scala 193:47]
  wire  _GEN_1151 = _T_3545 & _T_3572; // @[tlb.scala 193:47]
  wire  _GEN_1164 = _T_3545 & _T_3573; // @[tlb.scala 193:47]
  wire  _GEN_1177 = _T_3545 & _T_3574; // @[tlb.scala 193:47]
  wire  _GEN_1190 = _T_3545 & _T_3575; // @[tlb.scala 193:47]
  wire  _GEN_1203 = _T_3545 & _T_3576; // @[tlb.scala 193:47]
  wire  _GEN_1216 = _T_3545 & _T_3577; // @[tlb.scala 193:47]
  wire [31:0] _T_3578 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_0_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3579 = ~_T_3578; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1558 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_0_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3580 = _GEN_1558 & _T_3579; // @[tlb.scala 50:19]
  wire [31:0] _GEN_1559 = {{13'd0}, io_pport_entry_hi_vpn}; // @[tlb.scala 50:37]
  wire [31:0] _T_3582 = _GEN_1559 & _T_3579; // @[tlb.scala 50:37]
  wire  _T_3583 = _T_3580 == _T_3582; // @[tlb.scala 50:28]
  wire  _T_3584 = tlb_entries_asid_tlb_entry_ports_0_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3585 = tlb_entries_g_tlb_entry_ports_0_r_data | _T_3584; // @[tlb.scala 51:17]
  wire  _T_3586 = _T_3583 & _T_3585; // @[tlb.scala 50:46]
  wire [31:0] _T_3587 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_1_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3588 = ~_T_3587; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1560 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_1_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3589 = _GEN_1560 & _T_3588; // @[tlb.scala 50:19]
  wire [31:0] _T_3591 = _GEN_1559 & _T_3588; // @[tlb.scala 50:37]
  wire  _T_3592 = _T_3589 == _T_3591; // @[tlb.scala 50:28]
  wire  _T_3593 = tlb_entries_asid_tlb_entry_ports_1_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3594 = tlb_entries_g_tlb_entry_ports_1_r_data | _T_3593; // @[tlb.scala 51:17]
  wire  _T_3595 = _T_3592 & _T_3594; // @[tlb.scala 50:46]
  wire [31:0] _T_3596 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_2_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3597 = ~_T_3596; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1562 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_2_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3598 = _GEN_1562 & _T_3597; // @[tlb.scala 50:19]
  wire [31:0] _T_3600 = _GEN_1559 & _T_3597; // @[tlb.scala 50:37]
  wire  _T_3601 = _T_3598 == _T_3600; // @[tlb.scala 50:28]
  wire  _T_3602 = tlb_entries_asid_tlb_entry_ports_2_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3603 = tlb_entries_g_tlb_entry_ports_2_r_data | _T_3602; // @[tlb.scala 51:17]
  wire  _T_3604 = _T_3601 & _T_3603; // @[tlb.scala 50:46]
  wire [31:0] _T_3605 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_3_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3606 = ~_T_3605; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1564 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_3_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3607 = _GEN_1564 & _T_3606; // @[tlb.scala 50:19]
  wire [31:0] _T_3609 = _GEN_1559 & _T_3606; // @[tlb.scala 50:37]
  wire  _T_3610 = _T_3607 == _T_3609; // @[tlb.scala 50:28]
  wire  _T_3611 = tlb_entries_asid_tlb_entry_ports_3_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3612 = tlb_entries_g_tlb_entry_ports_3_r_data | _T_3611; // @[tlb.scala 51:17]
  wire  _T_3613 = _T_3610 & _T_3612; // @[tlb.scala 50:46]
  wire [31:0] _T_3614 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_4_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3615 = ~_T_3614; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1566 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_4_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3616 = _GEN_1566 & _T_3615; // @[tlb.scala 50:19]
  wire [31:0] _T_3618 = _GEN_1559 & _T_3615; // @[tlb.scala 50:37]
  wire  _T_3619 = _T_3616 == _T_3618; // @[tlb.scala 50:28]
  wire  _T_3620 = tlb_entries_asid_tlb_entry_ports_4_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3621 = tlb_entries_g_tlb_entry_ports_4_r_data | _T_3620; // @[tlb.scala 51:17]
  wire  _T_3622 = _T_3619 & _T_3621; // @[tlb.scala 50:46]
  wire [31:0] _T_3623 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_5_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3624 = ~_T_3623; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1568 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_5_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3625 = _GEN_1568 & _T_3624; // @[tlb.scala 50:19]
  wire [31:0] _T_3627 = _GEN_1559 & _T_3624; // @[tlb.scala 50:37]
  wire  _T_3628 = _T_3625 == _T_3627; // @[tlb.scala 50:28]
  wire  _T_3629 = tlb_entries_asid_tlb_entry_ports_5_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3630 = tlb_entries_g_tlb_entry_ports_5_r_data | _T_3629; // @[tlb.scala 51:17]
  wire  _T_3631 = _T_3628 & _T_3630; // @[tlb.scala 50:46]
  wire [31:0] _T_3632 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_6_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3633 = ~_T_3632; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1570 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_6_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3634 = _GEN_1570 & _T_3633; // @[tlb.scala 50:19]
  wire [31:0] _T_3636 = _GEN_1559 & _T_3633; // @[tlb.scala 50:37]
  wire  _T_3637 = _T_3634 == _T_3636; // @[tlb.scala 50:28]
  wire  _T_3638 = tlb_entries_asid_tlb_entry_ports_6_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3639 = tlb_entries_g_tlb_entry_ports_6_r_data | _T_3638; // @[tlb.scala 51:17]
  wire  _T_3640 = _T_3637 & _T_3639; // @[tlb.scala 50:46]
  wire [31:0] _T_3641 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_7_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3642 = ~_T_3641; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1572 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_7_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3643 = _GEN_1572 & _T_3642; // @[tlb.scala 50:19]
  wire [31:0] _T_3645 = _GEN_1559 & _T_3642; // @[tlb.scala 50:37]
  wire  _T_3646 = _T_3643 == _T_3645; // @[tlb.scala 50:28]
  wire  _T_3647 = tlb_entries_asid_tlb_entry_ports_7_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3648 = tlb_entries_g_tlb_entry_ports_7_r_data | _T_3647; // @[tlb.scala 51:17]
  wire  _T_3649 = _T_3646 & _T_3648; // @[tlb.scala 50:46]
  wire [31:0] _T_3650 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_8_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3651 = ~_T_3650; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1574 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_8_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3652 = _GEN_1574 & _T_3651; // @[tlb.scala 50:19]
  wire [31:0] _T_3654 = _GEN_1559 & _T_3651; // @[tlb.scala 50:37]
  wire  _T_3655 = _T_3652 == _T_3654; // @[tlb.scala 50:28]
  wire  _T_3656 = tlb_entries_asid_tlb_entry_ports_8_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3657 = tlb_entries_g_tlb_entry_ports_8_r_data | _T_3656; // @[tlb.scala 51:17]
  wire  _T_3658 = _T_3655 & _T_3657; // @[tlb.scala 50:46]
  wire [31:0] _T_3659 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_9_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3660 = ~_T_3659; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1576 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_9_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3661 = _GEN_1576 & _T_3660; // @[tlb.scala 50:19]
  wire [31:0] _T_3663 = _GEN_1559 & _T_3660; // @[tlb.scala 50:37]
  wire  _T_3664 = _T_3661 == _T_3663; // @[tlb.scala 50:28]
  wire  _T_3665 = tlb_entries_asid_tlb_entry_ports_9_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3666 = tlb_entries_g_tlb_entry_ports_9_r_data | _T_3665; // @[tlb.scala 51:17]
  wire  _T_3667 = _T_3664 & _T_3666; // @[tlb.scala 50:46]
  wire [31:0] _T_3668 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_10_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3669 = ~_T_3668; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1578 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_10_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3670 = _GEN_1578 & _T_3669; // @[tlb.scala 50:19]
  wire [31:0] _T_3672 = _GEN_1559 & _T_3669; // @[tlb.scala 50:37]
  wire  _T_3673 = _T_3670 == _T_3672; // @[tlb.scala 50:28]
  wire  _T_3674 = tlb_entries_asid_tlb_entry_ports_10_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3675 = tlb_entries_g_tlb_entry_ports_10_r_data | _T_3674; // @[tlb.scala 51:17]
  wire  _T_3676 = _T_3673 & _T_3675; // @[tlb.scala 50:46]
  wire [31:0] _T_3677 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_11_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3678 = ~_T_3677; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1580 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_11_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3679 = _GEN_1580 & _T_3678; // @[tlb.scala 50:19]
  wire [31:0] _T_3681 = _GEN_1559 & _T_3678; // @[tlb.scala 50:37]
  wire  _T_3682 = _T_3679 == _T_3681; // @[tlb.scala 50:28]
  wire  _T_3683 = tlb_entries_asid_tlb_entry_ports_11_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3684 = tlb_entries_g_tlb_entry_ports_11_r_data | _T_3683; // @[tlb.scala 51:17]
  wire  _T_3685 = _T_3682 & _T_3684; // @[tlb.scala 50:46]
  wire [31:0] _T_3686 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_12_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3687 = ~_T_3686; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1582 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_12_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3688 = _GEN_1582 & _T_3687; // @[tlb.scala 50:19]
  wire [31:0] _T_3690 = _GEN_1559 & _T_3687; // @[tlb.scala 50:37]
  wire  _T_3691 = _T_3688 == _T_3690; // @[tlb.scala 50:28]
  wire  _T_3692 = tlb_entries_asid_tlb_entry_ports_12_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3693 = tlb_entries_g_tlb_entry_ports_12_r_data | _T_3692; // @[tlb.scala 51:17]
  wire  _T_3694 = _T_3691 & _T_3693; // @[tlb.scala 50:46]
  wire [31:0] _T_3695 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_13_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3696 = ~_T_3695; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1584 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_13_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3697 = _GEN_1584 & _T_3696; // @[tlb.scala 50:19]
  wire [31:0] _T_3699 = _GEN_1559 & _T_3696; // @[tlb.scala 50:37]
  wire  _T_3700 = _T_3697 == _T_3699; // @[tlb.scala 50:28]
  wire  _T_3701 = tlb_entries_asid_tlb_entry_ports_13_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3702 = tlb_entries_g_tlb_entry_ports_13_r_data | _T_3701; // @[tlb.scala 51:17]
  wire  _T_3703 = _T_3700 & _T_3702; // @[tlb.scala 50:46]
  wire [31:0] _T_3704 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_14_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3705 = ~_T_3704; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1586 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_14_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3706 = _GEN_1586 & _T_3705; // @[tlb.scala 50:19]
  wire [31:0] _T_3708 = _GEN_1559 & _T_3705; // @[tlb.scala 50:37]
  wire  _T_3709 = _T_3706 == _T_3708; // @[tlb.scala 50:28]
  wire  _T_3710 = tlb_entries_asid_tlb_entry_ports_14_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3711 = tlb_entries_g_tlb_entry_ports_14_r_data | _T_3710; // @[tlb.scala 51:17]
  wire  _T_3712 = _T_3709 & _T_3711; // @[tlb.scala 50:46]
  wire [31:0] _T_3713 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_15_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3714 = ~_T_3713; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1588 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_15_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3715 = _GEN_1588 & _T_3714; // @[tlb.scala 50:19]
  wire [31:0] _T_3717 = _GEN_1559 & _T_3714; // @[tlb.scala 50:37]
  wire  _T_3718 = _T_3715 == _T_3717; // @[tlb.scala 50:28]
  wire  _T_3719 = tlb_entries_asid_tlb_entry_ports_15_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3720 = tlb_entries_g_tlb_entry_ports_15_r_data | _T_3719; // @[tlb.scala 51:17]
  wire  _T_3721 = _T_3718 & _T_3720; // @[tlb.scala 50:46]
  wire [31:0] _T_3722 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_16_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3723 = ~_T_3722; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1590 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_16_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3724 = _GEN_1590 & _T_3723; // @[tlb.scala 50:19]
  wire [31:0] _T_3726 = _GEN_1559 & _T_3723; // @[tlb.scala 50:37]
  wire  _T_3727 = _T_3724 == _T_3726; // @[tlb.scala 50:28]
  wire  _T_3728 = tlb_entries_asid_tlb_entry_ports_16_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3729 = tlb_entries_g_tlb_entry_ports_16_r_data | _T_3728; // @[tlb.scala 51:17]
  wire  _T_3730 = _T_3727 & _T_3729; // @[tlb.scala 50:46]
  wire [31:0] _T_3731 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_17_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3732 = ~_T_3731; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1592 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_17_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3733 = _GEN_1592 & _T_3732; // @[tlb.scala 50:19]
  wire [31:0] _T_3735 = _GEN_1559 & _T_3732; // @[tlb.scala 50:37]
  wire  _T_3736 = _T_3733 == _T_3735; // @[tlb.scala 50:28]
  wire  _T_3737 = tlb_entries_asid_tlb_entry_ports_17_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3738 = tlb_entries_g_tlb_entry_ports_17_r_data | _T_3737; // @[tlb.scala 51:17]
  wire  _T_3739 = _T_3736 & _T_3738; // @[tlb.scala 50:46]
  wire [31:0] _T_3740 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_18_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3741 = ~_T_3740; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1594 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_18_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3742 = _GEN_1594 & _T_3741; // @[tlb.scala 50:19]
  wire [31:0] _T_3744 = _GEN_1559 & _T_3741; // @[tlb.scala 50:37]
  wire  _T_3745 = _T_3742 == _T_3744; // @[tlb.scala 50:28]
  wire  _T_3746 = tlb_entries_asid_tlb_entry_ports_18_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3747 = tlb_entries_g_tlb_entry_ports_18_r_data | _T_3746; // @[tlb.scala 51:17]
  wire  _T_3748 = _T_3745 & _T_3747; // @[tlb.scala 50:46]
  wire [31:0] _T_3749 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_19_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3750 = ~_T_3749; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1596 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_19_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3751 = _GEN_1596 & _T_3750; // @[tlb.scala 50:19]
  wire [31:0] _T_3753 = _GEN_1559 & _T_3750; // @[tlb.scala 50:37]
  wire  _T_3754 = _T_3751 == _T_3753; // @[tlb.scala 50:28]
  wire  _T_3755 = tlb_entries_asid_tlb_entry_ports_19_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3756 = tlb_entries_g_tlb_entry_ports_19_r_data | _T_3755; // @[tlb.scala 51:17]
  wire  _T_3757 = _T_3754 & _T_3756; // @[tlb.scala 50:46]
  wire [31:0] _T_3758 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_20_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3759 = ~_T_3758; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1598 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_20_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3760 = _GEN_1598 & _T_3759; // @[tlb.scala 50:19]
  wire [31:0] _T_3762 = _GEN_1559 & _T_3759; // @[tlb.scala 50:37]
  wire  _T_3763 = _T_3760 == _T_3762; // @[tlb.scala 50:28]
  wire  _T_3764 = tlb_entries_asid_tlb_entry_ports_20_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3765 = tlb_entries_g_tlb_entry_ports_20_r_data | _T_3764; // @[tlb.scala 51:17]
  wire  _T_3766 = _T_3763 & _T_3765; // @[tlb.scala 50:46]
  wire [31:0] _T_3767 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_21_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3768 = ~_T_3767; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1600 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_21_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3769 = _GEN_1600 & _T_3768; // @[tlb.scala 50:19]
  wire [31:0] _T_3771 = _GEN_1559 & _T_3768; // @[tlb.scala 50:37]
  wire  _T_3772 = _T_3769 == _T_3771; // @[tlb.scala 50:28]
  wire  _T_3773 = tlb_entries_asid_tlb_entry_ports_21_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3774 = tlb_entries_g_tlb_entry_ports_21_r_data | _T_3773; // @[tlb.scala 51:17]
  wire  _T_3775 = _T_3772 & _T_3774; // @[tlb.scala 50:46]
  wire [31:0] _T_3776 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_22_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3777 = ~_T_3776; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1602 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_22_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3778 = _GEN_1602 & _T_3777; // @[tlb.scala 50:19]
  wire [31:0] _T_3780 = _GEN_1559 & _T_3777; // @[tlb.scala 50:37]
  wire  _T_3781 = _T_3778 == _T_3780; // @[tlb.scala 50:28]
  wire  _T_3782 = tlb_entries_asid_tlb_entry_ports_22_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3783 = tlb_entries_g_tlb_entry_ports_22_r_data | _T_3782; // @[tlb.scala 51:17]
  wire  _T_3784 = _T_3781 & _T_3783; // @[tlb.scala 50:46]
  wire [31:0] _T_3785 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_23_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3786 = ~_T_3785; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1604 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_23_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3787 = _GEN_1604 & _T_3786; // @[tlb.scala 50:19]
  wire [31:0] _T_3789 = _GEN_1559 & _T_3786; // @[tlb.scala 50:37]
  wire  _T_3790 = _T_3787 == _T_3789; // @[tlb.scala 50:28]
  wire  _T_3791 = tlb_entries_asid_tlb_entry_ports_23_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3792 = tlb_entries_g_tlb_entry_ports_23_r_data | _T_3791; // @[tlb.scala 51:17]
  wire  _T_3793 = _T_3790 & _T_3792; // @[tlb.scala 50:46]
  wire [31:0] _T_3794 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_24_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3795 = ~_T_3794; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1606 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_24_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3796 = _GEN_1606 & _T_3795; // @[tlb.scala 50:19]
  wire [31:0] _T_3798 = _GEN_1559 & _T_3795; // @[tlb.scala 50:37]
  wire  _T_3799 = _T_3796 == _T_3798; // @[tlb.scala 50:28]
  wire  _T_3800 = tlb_entries_asid_tlb_entry_ports_24_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3801 = tlb_entries_g_tlb_entry_ports_24_r_data | _T_3800; // @[tlb.scala 51:17]
  wire  _T_3802 = _T_3799 & _T_3801; // @[tlb.scala 50:46]
  wire [31:0] _T_3803 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_25_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3804 = ~_T_3803; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1608 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_25_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3805 = _GEN_1608 & _T_3804; // @[tlb.scala 50:19]
  wire [31:0] _T_3807 = _GEN_1559 & _T_3804; // @[tlb.scala 50:37]
  wire  _T_3808 = _T_3805 == _T_3807; // @[tlb.scala 50:28]
  wire  _T_3809 = tlb_entries_asid_tlb_entry_ports_25_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3810 = tlb_entries_g_tlb_entry_ports_25_r_data | _T_3809; // @[tlb.scala 51:17]
  wire  _T_3811 = _T_3808 & _T_3810; // @[tlb.scala 50:46]
  wire [31:0] _T_3812 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_26_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3813 = ~_T_3812; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1610 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_26_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3814 = _GEN_1610 & _T_3813; // @[tlb.scala 50:19]
  wire [31:0] _T_3816 = _GEN_1559 & _T_3813; // @[tlb.scala 50:37]
  wire  _T_3817 = _T_3814 == _T_3816; // @[tlb.scala 50:28]
  wire  _T_3818 = tlb_entries_asid_tlb_entry_ports_26_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3819 = tlb_entries_g_tlb_entry_ports_26_r_data | _T_3818; // @[tlb.scala 51:17]
  wire  _T_3820 = _T_3817 & _T_3819; // @[tlb.scala 50:46]
  wire [31:0] _T_3821 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_27_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3822 = ~_T_3821; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1612 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_27_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3823 = _GEN_1612 & _T_3822; // @[tlb.scala 50:19]
  wire [31:0] _T_3825 = _GEN_1559 & _T_3822; // @[tlb.scala 50:37]
  wire  _T_3826 = _T_3823 == _T_3825; // @[tlb.scala 50:28]
  wire  _T_3827 = tlb_entries_asid_tlb_entry_ports_27_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3828 = tlb_entries_g_tlb_entry_ports_27_r_data | _T_3827; // @[tlb.scala 51:17]
  wire  _T_3829 = _T_3826 & _T_3828; // @[tlb.scala 50:46]
  wire [31:0] _T_3830 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_28_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3831 = ~_T_3830; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1614 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_28_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3832 = _GEN_1614 & _T_3831; // @[tlb.scala 50:19]
  wire [31:0] _T_3834 = _GEN_1559 & _T_3831; // @[tlb.scala 50:37]
  wire  _T_3835 = _T_3832 == _T_3834; // @[tlb.scala 50:28]
  wire  _T_3836 = tlb_entries_asid_tlb_entry_ports_28_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3837 = tlb_entries_g_tlb_entry_ports_28_r_data | _T_3836; // @[tlb.scala 51:17]
  wire  _T_3838 = _T_3835 & _T_3837; // @[tlb.scala 50:46]
  wire [31:0] _T_3839 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_29_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3840 = ~_T_3839; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1616 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_29_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3841 = _GEN_1616 & _T_3840; // @[tlb.scala 50:19]
  wire [31:0] _T_3843 = _GEN_1559 & _T_3840; // @[tlb.scala 50:37]
  wire  _T_3844 = _T_3841 == _T_3843; // @[tlb.scala 50:28]
  wire  _T_3845 = tlb_entries_asid_tlb_entry_ports_29_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3846 = tlb_entries_g_tlb_entry_ports_29_r_data | _T_3845; // @[tlb.scala 51:17]
  wire  _T_3847 = _T_3844 & _T_3846; // @[tlb.scala 50:46]
  wire [31:0] _T_3848 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_30_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3849 = ~_T_3848; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1618 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_30_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3850 = _GEN_1618 & _T_3849; // @[tlb.scala 50:19]
  wire [31:0] _T_3852 = _GEN_1559 & _T_3849; // @[tlb.scala 50:37]
  wire  _T_3853 = _T_3850 == _T_3852; // @[tlb.scala 50:28]
  wire  _T_3854 = tlb_entries_asid_tlb_entry_ports_30_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3855 = tlb_entries_g_tlb_entry_ports_30_r_data | _T_3854; // @[tlb.scala 51:17]
  wire  _T_3856 = _T_3853 & _T_3855; // @[tlb.scala 50:46]
  wire [31:0] _T_3857 = {{16'd0}, tlb_entries_pagemask_tlb_entry_ports_31_r_data}; // @[tlb.scala 49:42 tlb.scala 49:42]
  wire [31:0] _T_3858 = ~_T_3857; // @[tlb.scala 50:21]
  wire [31:0] _GEN_1620 = {{13'd0}, tlb_entries_vpn_tlb_entry_ports_31_r_data}; // @[tlb.scala 50:19]
  wire [31:0] _T_3859 = _GEN_1620 & _T_3858; // @[tlb.scala 50:19]
  wire [31:0] _T_3861 = _GEN_1559 & _T_3858; // @[tlb.scala 50:37]
  wire  _T_3862 = _T_3859 == _T_3861; // @[tlb.scala 50:28]
  wire  _T_3863 = tlb_entries_asid_tlb_entry_ports_31_r_data == io_pport_entry_hi_asid; // @[tlb.scala 51:34]
  wire  _T_3864 = tlb_entries_g_tlb_entry_ports_31_r_data | _T_3863; // @[tlb.scala 51:17]
  wire  _T_3865 = _T_3862 & _T_3864; // @[tlb.scala 50:46]
  wire [7:0] _T_3872 = {_T_3802,_T_3811,_T_3820,_T_3829,_T_3838,_T_3847,_T_3856,_T_3865}; // @[Cat.scala 29:58]
  wire [15:0] _T_3880 = {_T_3730,_T_3739,_T_3748,_T_3757,_T_3766,_T_3775,_T_3784,_T_3793,_T_3872}; // @[Cat.scala 29:58]
  wire [7:0] _T_3887 = {_T_3658,_T_3667,_T_3676,_T_3685,_T_3694,_T_3703,_T_3712,_T_3721}; // @[Cat.scala 29:58]
  wire [31:0] _T_3896 = {_T_3586,_T_3595,_T_3604,_T_3613,_T_3622,_T_3631,_T_3640,_T_3649,_T_3887,_T_3880}; // @[Cat.scala 29:58]
  wire [31:0] _T_3900 = {{16'd0}, _T_3896[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3902 = {_T_3896[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_3904 = _T_3902 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_3905 = _T_3900 | _T_3904; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1622 = {{8'd0}, _T_3905[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3910 = _GEN_1622 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3912 = {_T_3905[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_3914 = _T_3912 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_3915 = _T_3910 | _T_3914; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1623 = {{4'd0}, _T_3915[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3920 = _GEN_1623 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3922 = {_T_3915[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_3924 = _T_3922 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_3925 = _T_3920 | _T_3924; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1624 = {{2'd0}, _T_3925[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3930 = _GEN_1624 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3932 = {_T_3925[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_3934 = _T_3932 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_3935 = _T_3930 | _T_3934; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1625 = {{1'd0}, _T_3935[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3940 = _GEN_1625 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_3942 = {_T_3935[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_3944 = _T_3942 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] matches_ = _T_3940 | _T_3944; // @[Bitwise.scala 103:39]
  wire  _T_3945 = matches_ != 32'h0; // @[tlb.scala 203:32]
  wire [1:0] _T_3981 = matches_[2] ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_3982 = matches_[3] ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_3983 = matches_[4] ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_3984 = matches_[5] ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_3985 = matches_[6] ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_3986 = matches_[7] ? 3'h7 : 3'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3987 = matches_[8] ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3988 = matches_[9] ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3989 = matches_[10] ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3990 = matches_[11] ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3991 = matches_[12] ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3992 = matches_[13] ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3993 = matches_[14] ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_3994 = matches_[15] ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3995 = matches_[16] ? 5'h10 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3996 = matches_[17] ? 5'h11 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3997 = matches_[18] ? 5'h12 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3998 = matches_[19] ? 5'h13 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_3999 = matches_[20] ? 5'h14 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4000 = matches_[21] ? 5'h15 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4001 = matches_[22] ? 5'h16 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4002 = matches_[23] ? 5'h17 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4003 = matches_[24] ? 5'h18 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4004 = matches_[25] ? 5'h19 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4005 = matches_[26] ? 5'h1a : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4006 = matches_[27] ? 5'h1b : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4007 = matches_[28] ? 5'h1c : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4008 = matches_[29] ? 5'h1d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4009 = matches_[30] ? 5'h1e : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_4010 = matches_[31] ? 5'h1f : 5'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_1626 = {{1'd0}, matches_[1]}; // @[Mux.scala 27:72]
  wire [1:0] _T_4012 = _GEN_1626 | _T_3981; // @[Mux.scala 27:72]
  wire [1:0] _T_4013 = _T_4012 | _T_3982; // @[Mux.scala 27:72]
  wire [2:0] _GEN_1627 = {{1'd0}, _T_4013}; // @[Mux.scala 27:72]
  wire [2:0] _T_4014 = _GEN_1627 | _T_3983; // @[Mux.scala 27:72]
  wire [2:0] _T_4015 = _T_4014 | _T_3984; // @[Mux.scala 27:72]
  wire [2:0] _T_4016 = _T_4015 | _T_3985; // @[Mux.scala 27:72]
  wire [2:0] _T_4017 = _T_4016 | _T_3986; // @[Mux.scala 27:72]
  wire [3:0] _GEN_1628 = {{1'd0}, _T_4017}; // @[Mux.scala 27:72]
  wire [3:0] _T_4018 = _GEN_1628 | _T_3987; // @[Mux.scala 27:72]
  wire [3:0] _T_4019 = _T_4018 | _T_3988; // @[Mux.scala 27:72]
  wire [3:0] _T_4020 = _T_4019 | _T_3989; // @[Mux.scala 27:72]
  wire [3:0] _T_4021 = _T_4020 | _T_3990; // @[Mux.scala 27:72]
  wire [3:0] _T_4022 = _T_4021 | _T_3991; // @[Mux.scala 27:72]
  wire [3:0] _T_4023 = _T_4022 | _T_3992; // @[Mux.scala 27:72]
  wire [3:0] _T_4024 = _T_4023 | _T_3993; // @[Mux.scala 27:72]
  wire [3:0] _T_4025 = _T_4024 | _T_3994; // @[Mux.scala 27:72]
  wire [4:0] _GEN_1629 = {{1'd0}, _T_4025}; // @[Mux.scala 27:72]
  wire [4:0] _T_4026 = _GEN_1629 | _T_3995; // @[Mux.scala 27:72]
  wire [4:0] _T_4027 = _T_4026 | _T_3996; // @[Mux.scala 27:72]
  wire [4:0] _T_4028 = _T_4027 | _T_3997; // @[Mux.scala 27:72]
  wire [4:0] _T_4029 = _T_4028 | _T_3998; // @[Mux.scala 27:72]
  wire [4:0] _T_4030 = _T_4029 | _T_3999; // @[Mux.scala 27:72]
  wire [4:0] _T_4031 = _T_4030 | _T_4000; // @[Mux.scala 27:72]
  wire [4:0] _T_4032 = _T_4031 | _T_4001; // @[Mux.scala 27:72]
  wire [4:0] _T_4033 = _T_4032 | _T_4002; // @[Mux.scala 27:72]
  wire [4:0] _T_4034 = _T_4033 | _T_4003; // @[Mux.scala 27:72]
  wire [4:0] _T_4035 = _T_4034 | _T_4004; // @[Mux.scala 27:72]
  wire [4:0] _T_4036 = _T_4035 | _T_4005; // @[Mux.scala 27:72]
  wire [4:0] _T_4037 = _T_4036 | _T_4006; // @[Mux.scala 27:72]
  wire [4:0] _T_4038 = _T_4037 | _T_4007; // @[Mux.scala 27:72]
  wire [4:0] _T_4039 = _T_4038 | _T_4008; // @[Mux.scala 27:72]
  wire [4:0] _T_4040 = _T_4039 | _T_4009; // @[Mux.scala 27:72]
  assign tlb_entries_pagemask__T_5_addr = 5'h0;
  assign tlb_entries_pagemask__T_5_data = tlb_entries_pagemask[tlb_entries_pagemask__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_6_addr = 5'h1;
  assign tlb_entries_pagemask__T_6_data = tlb_entries_pagemask[tlb_entries_pagemask__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_7_addr = 5'h2;
  assign tlb_entries_pagemask__T_7_data = tlb_entries_pagemask[tlb_entries_pagemask__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_8_addr = 5'h3;
  assign tlb_entries_pagemask__T_8_data = tlb_entries_pagemask[tlb_entries_pagemask__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_9_addr = 5'h4;
  assign tlb_entries_pagemask__T_9_data = tlb_entries_pagemask[tlb_entries_pagemask__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_10_addr = 5'h5;
  assign tlb_entries_pagemask__T_10_data = tlb_entries_pagemask[tlb_entries_pagemask__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_11_addr = 5'h6;
  assign tlb_entries_pagemask__T_11_data = tlb_entries_pagemask[tlb_entries_pagemask__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_12_addr = 5'h7;
  assign tlb_entries_pagemask__T_12_data = tlb_entries_pagemask[tlb_entries_pagemask__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_13_addr = 5'h8;
  assign tlb_entries_pagemask__T_13_data = tlb_entries_pagemask[tlb_entries_pagemask__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_14_addr = 5'h9;
  assign tlb_entries_pagemask__T_14_data = tlb_entries_pagemask[tlb_entries_pagemask__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_15_addr = 5'ha;
  assign tlb_entries_pagemask__T_15_data = tlb_entries_pagemask[tlb_entries_pagemask__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_16_addr = 5'hb;
  assign tlb_entries_pagemask__T_16_data = tlb_entries_pagemask[tlb_entries_pagemask__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_17_addr = 5'hc;
  assign tlb_entries_pagemask__T_17_data = tlb_entries_pagemask[tlb_entries_pagemask__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_18_addr = 5'hd;
  assign tlb_entries_pagemask__T_18_data = tlb_entries_pagemask[tlb_entries_pagemask__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_19_addr = 5'he;
  assign tlb_entries_pagemask__T_19_data = tlb_entries_pagemask[tlb_entries_pagemask__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_20_addr = 5'hf;
  assign tlb_entries_pagemask__T_20_data = tlb_entries_pagemask[tlb_entries_pagemask__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_21_addr = 5'h10;
  assign tlb_entries_pagemask__T_21_data = tlb_entries_pagemask[tlb_entries_pagemask__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_22_addr = 5'h11;
  assign tlb_entries_pagemask__T_22_data = tlb_entries_pagemask[tlb_entries_pagemask__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_23_addr = 5'h12;
  assign tlb_entries_pagemask__T_23_data = tlb_entries_pagemask[tlb_entries_pagemask__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_24_addr = 5'h13;
  assign tlb_entries_pagemask__T_24_data = tlb_entries_pagemask[tlb_entries_pagemask__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_25_addr = 5'h14;
  assign tlb_entries_pagemask__T_25_data = tlb_entries_pagemask[tlb_entries_pagemask__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_26_addr = 5'h15;
  assign tlb_entries_pagemask__T_26_data = tlb_entries_pagemask[tlb_entries_pagemask__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_27_addr = 5'h16;
  assign tlb_entries_pagemask__T_27_data = tlb_entries_pagemask[tlb_entries_pagemask__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_28_addr = 5'h17;
  assign tlb_entries_pagemask__T_28_data = tlb_entries_pagemask[tlb_entries_pagemask__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_29_addr = 5'h18;
  assign tlb_entries_pagemask__T_29_data = tlb_entries_pagemask[tlb_entries_pagemask__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_30_addr = 5'h19;
  assign tlb_entries_pagemask__T_30_data = tlb_entries_pagemask[tlb_entries_pagemask__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_31_addr = 5'h1a;
  assign tlb_entries_pagemask__T_31_data = tlb_entries_pagemask[tlb_entries_pagemask__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_32_addr = 5'h1b;
  assign tlb_entries_pagemask__T_32_data = tlb_entries_pagemask[tlb_entries_pagemask__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_33_addr = 5'h1c;
  assign tlb_entries_pagemask__T_33_data = tlb_entries_pagemask[tlb_entries_pagemask__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_34_addr = 5'h1d;
  assign tlb_entries_pagemask__T_34_data = tlb_entries_pagemask[tlb_entries_pagemask__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_35_addr = 5'h1e;
  assign tlb_entries_pagemask__T_35_data = tlb_entries_pagemask[tlb_entries_pagemask__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_36_addr = 5'h1f;
  assign tlb_entries_pagemask__T_36_data = tlb_entries_pagemask[tlb_entries_pagemask__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1546_addr = 5'h0;
  assign tlb_entries_pagemask__T_1546_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1547_addr = 5'h1;
  assign tlb_entries_pagemask__T_1547_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1548_addr = 5'h2;
  assign tlb_entries_pagemask__T_1548_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1549_addr = 5'h3;
  assign tlb_entries_pagemask__T_1549_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1550_addr = 5'h4;
  assign tlb_entries_pagemask__T_1550_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1551_addr = 5'h5;
  assign tlb_entries_pagemask__T_1551_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1552_addr = 5'h6;
  assign tlb_entries_pagemask__T_1552_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1553_addr = 5'h7;
  assign tlb_entries_pagemask__T_1553_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1554_addr = 5'h8;
  assign tlb_entries_pagemask__T_1554_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1555_addr = 5'h9;
  assign tlb_entries_pagemask__T_1555_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1556_addr = 5'ha;
  assign tlb_entries_pagemask__T_1556_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1557_addr = 5'hb;
  assign tlb_entries_pagemask__T_1557_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1558_addr = 5'hc;
  assign tlb_entries_pagemask__T_1558_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1559_addr = 5'hd;
  assign tlb_entries_pagemask__T_1559_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1560_addr = 5'he;
  assign tlb_entries_pagemask__T_1560_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1561_addr = 5'hf;
  assign tlb_entries_pagemask__T_1561_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1562_addr = 5'h10;
  assign tlb_entries_pagemask__T_1562_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1563_addr = 5'h11;
  assign tlb_entries_pagemask__T_1563_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1564_addr = 5'h12;
  assign tlb_entries_pagemask__T_1564_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1565_addr = 5'h13;
  assign tlb_entries_pagemask__T_1565_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1566_addr = 5'h14;
  assign tlb_entries_pagemask__T_1566_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1567_addr = 5'h15;
  assign tlb_entries_pagemask__T_1567_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1568_addr = 5'h16;
  assign tlb_entries_pagemask__T_1568_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1569_addr = 5'h17;
  assign tlb_entries_pagemask__T_1569_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1570_addr = 5'h18;
  assign tlb_entries_pagemask__T_1570_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1571_addr = 5'h19;
  assign tlb_entries_pagemask__T_1571_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1572_addr = 5'h1a;
  assign tlb_entries_pagemask__T_1572_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1573_addr = 5'h1b;
  assign tlb_entries_pagemask__T_1573_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1574_addr = 5'h1c;
  assign tlb_entries_pagemask__T_1574_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1575_addr = 5'h1d;
  assign tlb_entries_pagemask__T_1575_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1576_addr = 5'h1e;
  assign tlb_entries_pagemask__T_1576_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask__T_1577_addr = 5'h1f;
  assign tlb_entries_pagemask__T_1577_data = tlb_entries_pagemask[tlb_entries_pagemask__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_pagemask_tlb_entry_ports_0_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_pagemask_tlb_entry_ports_1_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_pagemask_tlb_entry_ports_2_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_pagemask_tlb_entry_ports_3_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_pagemask_tlb_entry_ports_4_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_pagemask_tlb_entry_ports_5_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_pagemask_tlb_entry_ports_6_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_pagemask_tlb_entry_ports_7_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_pagemask_tlb_entry_ports_8_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_pagemask_tlb_entry_ports_9_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_pagemask_tlb_entry_ports_10_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_pagemask_tlb_entry_ports_11_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_pagemask_tlb_entry_ports_12_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_pagemask_tlb_entry_ports_13_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_pagemask_tlb_entry_ports_14_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_pagemask_tlb_entry_ports_15_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_pagemask_tlb_entry_ports_16_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_pagemask_tlb_entry_ports_17_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_pagemask_tlb_entry_ports_18_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_pagemask_tlb_entry_ports_19_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_pagemask_tlb_entry_ports_20_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_pagemask_tlb_entry_ports_21_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_pagemask_tlb_entry_ports_22_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_pagemask_tlb_entry_ports_23_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_pagemask_tlb_entry_ports_24_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_pagemask_tlb_entry_ports_25_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_pagemask_tlb_entry_ports_26_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_pagemask_tlb_entry_ports_27_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_pagemask_tlb_entry_ports_28_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_pagemask_tlb_entry_ports_29_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_pagemask_tlb_entry_ports_30_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_pagemask_tlb_entry_ports_31_r_data = tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_pagemask_tlb_entry_ports_0_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_pagemask_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_pagemask_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_pagemask_tlb_entry_ports_1_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_pagemask_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_pagemask_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_pagemask_tlb_entry_ports_2_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_pagemask_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_pagemask_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_pagemask_tlb_entry_ports_3_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_pagemask_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_pagemask_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_pagemask_tlb_entry_ports_4_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_pagemask_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_pagemask_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_pagemask_tlb_entry_ports_5_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_pagemask_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_pagemask_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_pagemask_tlb_entry_ports_6_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_pagemask_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_pagemask_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_pagemask_tlb_entry_ports_7_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_pagemask_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_pagemask_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_pagemask_tlb_entry_ports_8_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_pagemask_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_pagemask_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_pagemask_tlb_entry_ports_9_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_pagemask_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_pagemask_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_pagemask_tlb_entry_ports_10_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_pagemask_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_pagemask_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_pagemask_tlb_entry_ports_11_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_pagemask_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_pagemask_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_pagemask_tlb_entry_ports_12_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_pagemask_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_pagemask_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_pagemask_tlb_entry_ports_13_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_pagemask_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_pagemask_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_pagemask_tlb_entry_ports_14_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_pagemask_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_pagemask_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_pagemask_tlb_entry_ports_15_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_pagemask_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_pagemask_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_pagemask_tlb_entry_ports_16_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_pagemask_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_pagemask_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_pagemask_tlb_entry_ports_17_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_pagemask_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_pagemask_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_pagemask_tlb_entry_ports_18_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_pagemask_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_pagemask_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_pagemask_tlb_entry_ports_19_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_pagemask_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_pagemask_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_pagemask_tlb_entry_ports_20_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_pagemask_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_pagemask_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_pagemask_tlb_entry_ports_21_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_pagemask_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_pagemask_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_pagemask_tlb_entry_ports_22_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_pagemask_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_pagemask_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_pagemask_tlb_entry_ports_23_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_pagemask_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_pagemask_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_pagemask_tlb_entry_ports_24_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_pagemask_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_pagemask_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_pagemask_tlb_entry_ports_25_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_pagemask_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_pagemask_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_pagemask_tlb_entry_ports_26_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_pagemask_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_pagemask_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_pagemask_tlb_entry_ports_27_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_pagemask_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_pagemask_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_pagemask_tlb_entry_ports_28_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_pagemask_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_pagemask_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_pagemask_tlb_entry_ports_29_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_pagemask_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_pagemask_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_pagemask_tlb_entry_ports_30_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_pagemask_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_pagemask_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_pagemask_tlb_entry_ports_31_w_data = io_wport_bits_entry_pagemask;
  assign tlb_entries_pagemask_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_pagemask_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_pagemask_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_vpn__T_5_addr = 5'h0;
  assign tlb_entries_vpn__T_5_data = tlb_entries_vpn[tlb_entries_vpn__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_6_addr = 5'h1;
  assign tlb_entries_vpn__T_6_data = tlb_entries_vpn[tlb_entries_vpn__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_7_addr = 5'h2;
  assign tlb_entries_vpn__T_7_data = tlb_entries_vpn[tlb_entries_vpn__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_8_addr = 5'h3;
  assign tlb_entries_vpn__T_8_data = tlb_entries_vpn[tlb_entries_vpn__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_9_addr = 5'h4;
  assign tlb_entries_vpn__T_9_data = tlb_entries_vpn[tlb_entries_vpn__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_10_addr = 5'h5;
  assign tlb_entries_vpn__T_10_data = tlb_entries_vpn[tlb_entries_vpn__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_11_addr = 5'h6;
  assign tlb_entries_vpn__T_11_data = tlb_entries_vpn[tlb_entries_vpn__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_12_addr = 5'h7;
  assign tlb_entries_vpn__T_12_data = tlb_entries_vpn[tlb_entries_vpn__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_13_addr = 5'h8;
  assign tlb_entries_vpn__T_13_data = tlb_entries_vpn[tlb_entries_vpn__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_14_addr = 5'h9;
  assign tlb_entries_vpn__T_14_data = tlb_entries_vpn[tlb_entries_vpn__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_15_addr = 5'ha;
  assign tlb_entries_vpn__T_15_data = tlb_entries_vpn[tlb_entries_vpn__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_16_addr = 5'hb;
  assign tlb_entries_vpn__T_16_data = tlb_entries_vpn[tlb_entries_vpn__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_17_addr = 5'hc;
  assign tlb_entries_vpn__T_17_data = tlb_entries_vpn[tlb_entries_vpn__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_18_addr = 5'hd;
  assign tlb_entries_vpn__T_18_data = tlb_entries_vpn[tlb_entries_vpn__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_19_addr = 5'he;
  assign tlb_entries_vpn__T_19_data = tlb_entries_vpn[tlb_entries_vpn__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_20_addr = 5'hf;
  assign tlb_entries_vpn__T_20_data = tlb_entries_vpn[tlb_entries_vpn__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_21_addr = 5'h10;
  assign tlb_entries_vpn__T_21_data = tlb_entries_vpn[tlb_entries_vpn__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_22_addr = 5'h11;
  assign tlb_entries_vpn__T_22_data = tlb_entries_vpn[tlb_entries_vpn__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_23_addr = 5'h12;
  assign tlb_entries_vpn__T_23_data = tlb_entries_vpn[tlb_entries_vpn__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_24_addr = 5'h13;
  assign tlb_entries_vpn__T_24_data = tlb_entries_vpn[tlb_entries_vpn__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_25_addr = 5'h14;
  assign tlb_entries_vpn__T_25_data = tlb_entries_vpn[tlb_entries_vpn__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_26_addr = 5'h15;
  assign tlb_entries_vpn__T_26_data = tlb_entries_vpn[tlb_entries_vpn__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_27_addr = 5'h16;
  assign tlb_entries_vpn__T_27_data = tlb_entries_vpn[tlb_entries_vpn__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_28_addr = 5'h17;
  assign tlb_entries_vpn__T_28_data = tlb_entries_vpn[tlb_entries_vpn__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_29_addr = 5'h18;
  assign tlb_entries_vpn__T_29_data = tlb_entries_vpn[tlb_entries_vpn__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_30_addr = 5'h19;
  assign tlb_entries_vpn__T_30_data = tlb_entries_vpn[tlb_entries_vpn__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_31_addr = 5'h1a;
  assign tlb_entries_vpn__T_31_data = tlb_entries_vpn[tlb_entries_vpn__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_32_addr = 5'h1b;
  assign tlb_entries_vpn__T_32_data = tlb_entries_vpn[tlb_entries_vpn__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_33_addr = 5'h1c;
  assign tlb_entries_vpn__T_33_data = tlb_entries_vpn[tlb_entries_vpn__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_34_addr = 5'h1d;
  assign tlb_entries_vpn__T_34_data = tlb_entries_vpn[tlb_entries_vpn__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_35_addr = 5'h1e;
  assign tlb_entries_vpn__T_35_data = tlb_entries_vpn[tlb_entries_vpn__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_36_addr = 5'h1f;
  assign tlb_entries_vpn__T_36_data = tlb_entries_vpn[tlb_entries_vpn__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1546_addr = 5'h0;
  assign tlb_entries_vpn__T_1546_data = tlb_entries_vpn[tlb_entries_vpn__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1547_addr = 5'h1;
  assign tlb_entries_vpn__T_1547_data = tlb_entries_vpn[tlb_entries_vpn__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1548_addr = 5'h2;
  assign tlb_entries_vpn__T_1548_data = tlb_entries_vpn[tlb_entries_vpn__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1549_addr = 5'h3;
  assign tlb_entries_vpn__T_1549_data = tlb_entries_vpn[tlb_entries_vpn__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1550_addr = 5'h4;
  assign tlb_entries_vpn__T_1550_data = tlb_entries_vpn[tlb_entries_vpn__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1551_addr = 5'h5;
  assign tlb_entries_vpn__T_1551_data = tlb_entries_vpn[tlb_entries_vpn__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1552_addr = 5'h6;
  assign tlb_entries_vpn__T_1552_data = tlb_entries_vpn[tlb_entries_vpn__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1553_addr = 5'h7;
  assign tlb_entries_vpn__T_1553_data = tlb_entries_vpn[tlb_entries_vpn__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1554_addr = 5'h8;
  assign tlb_entries_vpn__T_1554_data = tlb_entries_vpn[tlb_entries_vpn__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1555_addr = 5'h9;
  assign tlb_entries_vpn__T_1555_data = tlb_entries_vpn[tlb_entries_vpn__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1556_addr = 5'ha;
  assign tlb_entries_vpn__T_1556_data = tlb_entries_vpn[tlb_entries_vpn__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1557_addr = 5'hb;
  assign tlb_entries_vpn__T_1557_data = tlb_entries_vpn[tlb_entries_vpn__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1558_addr = 5'hc;
  assign tlb_entries_vpn__T_1558_data = tlb_entries_vpn[tlb_entries_vpn__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1559_addr = 5'hd;
  assign tlb_entries_vpn__T_1559_data = tlb_entries_vpn[tlb_entries_vpn__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1560_addr = 5'he;
  assign tlb_entries_vpn__T_1560_data = tlb_entries_vpn[tlb_entries_vpn__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1561_addr = 5'hf;
  assign tlb_entries_vpn__T_1561_data = tlb_entries_vpn[tlb_entries_vpn__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1562_addr = 5'h10;
  assign tlb_entries_vpn__T_1562_data = tlb_entries_vpn[tlb_entries_vpn__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1563_addr = 5'h11;
  assign tlb_entries_vpn__T_1563_data = tlb_entries_vpn[tlb_entries_vpn__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1564_addr = 5'h12;
  assign tlb_entries_vpn__T_1564_data = tlb_entries_vpn[tlb_entries_vpn__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1565_addr = 5'h13;
  assign tlb_entries_vpn__T_1565_data = tlb_entries_vpn[tlb_entries_vpn__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1566_addr = 5'h14;
  assign tlb_entries_vpn__T_1566_data = tlb_entries_vpn[tlb_entries_vpn__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1567_addr = 5'h15;
  assign tlb_entries_vpn__T_1567_data = tlb_entries_vpn[tlb_entries_vpn__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1568_addr = 5'h16;
  assign tlb_entries_vpn__T_1568_data = tlb_entries_vpn[tlb_entries_vpn__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1569_addr = 5'h17;
  assign tlb_entries_vpn__T_1569_data = tlb_entries_vpn[tlb_entries_vpn__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1570_addr = 5'h18;
  assign tlb_entries_vpn__T_1570_data = tlb_entries_vpn[tlb_entries_vpn__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1571_addr = 5'h19;
  assign tlb_entries_vpn__T_1571_data = tlb_entries_vpn[tlb_entries_vpn__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1572_addr = 5'h1a;
  assign tlb_entries_vpn__T_1572_data = tlb_entries_vpn[tlb_entries_vpn__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1573_addr = 5'h1b;
  assign tlb_entries_vpn__T_1573_data = tlb_entries_vpn[tlb_entries_vpn__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1574_addr = 5'h1c;
  assign tlb_entries_vpn__T_1574_data = tlb_entries_vpn[tlb_entries_vpn__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1575_addr = 5'h1d;
  assign tlb_entries_vpn__T_1575_data = tlb_entries_vpn[tlb_entries_vpn__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1576_addr = 5'h1e;
  assign tlb_entries_vpn__T_1576_data = tlb_entries_vpn[tlb_entries_vpn__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn__T_1577_addr = 5'h1f;
  assign tlb_entries_vpn__T_1577_data = tlb_entries_vpn[tlb_entries_vpn__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_vpn_tlb_entry_ports_0_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_vpn_tlb_entry_ports_1_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_vpn_tlb_entry_ports_2_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_vpn_tlb_entry_ports_3_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_vpn_tlb_entry_ports_4_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_vpn_tlb_entry_ports_5_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_vpn_tlb_entry_ports_6_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_vpn_tlb_entry_ports_7_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_vpn_tlb_entry_ports_8_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_vpn_tlb_entry_ports_9_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_vpn_tlb_entry_ports_10_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_vpn_tlb_entry_ports_11_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_vpn_tlb_entry_ports_12_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_vpn_tlb_entry_ports_13_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_vpn_tlb_entry_ports_14_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_vpn_tlb_entry_ports_15_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_vpn_tlb_entry_ports_16_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_vpn_tlb_entry_ports_17_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_vpn_tlb_entry_ports_18_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_vpn_tlb_entry_ports_19_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_vpn_tlb_entry_ports_20_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_vpn_tlb_entry_ports_21_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_vpn_tlb_entry_ports_22_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_vpn_tlb_entry_ports_23_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_vpn_tlb_entry_ports_24_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_vpn_tlb_entry_ports_25_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_vpn_tlb_entry_ports_26_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_vpn_tlb_entry_ports_27_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_vpn_tlb_entry_ports_28_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_vpn_tlb_entry_ports_29_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_vpn_tlb_entry_ports_30_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_vpn_tlb_entry_ports_31_r_data = tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_vpn_tlb_entry_ports_0_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_vpn_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_vpn_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_vpn_tlb_entry_ports_1_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_vpn_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_vpn_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_vpn_tlb_entry_ports_2_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_vpn_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_vpn_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_vpn_tlb_entry_ports_3_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_vpn_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_vpn_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_vpn_tlb_entry_ports_4_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_vpn_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_vpn_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_vpn_tlb_entry_ports_5_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_vpn_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_vpn_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_vpn_tlb_entry_ports_6_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_vpn_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_vpn_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_vpn_tlb_entry_ports_7_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_vpn_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_vpn_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_vpn_tlb_entry_ports_8_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_vpn_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_vpn_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_vpn_tlb_entry_ports_9_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_vpn_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_vpn_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_vpn_tlb_entry_ports_10_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_vpn_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_vpn_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_vpn_tlb_entry_ports_11_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_vpn_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_vpn_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_vpn_tlb_entry_ports_12_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_vpn_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_vpn_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_vpn_tlb_entry_ports_13_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_vpn_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_vpn_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_vpn_tlb_entry_ports_14_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_vpn_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_vpn_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_vpn_tlb_entry_ports_15_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_vpn_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_vpn_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_vpn_tlb_entry_ports_16_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_vpn_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_vpn_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_vpn_tlb_entry_ports_17_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_vpn_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_vpn_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_vpn_tlb_entry_ports_18_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_vpn_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_vpn_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_vpn_tlb_entry_ports_19_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_vpn_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_vpn_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_vpn_tlb_entry_ports_20_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_vpn_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_vpn_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_vpn_tlb_entry_ports_21_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_vpn_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_vpn_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_vpn_tlb_entry_ports_22_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_vpn_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_vpn_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_vpn_tlb_entry_ports_23_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_vpn_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_vpn_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_vpn_tlb_entry_ports_24_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_vpn_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_vpn_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_vpn_tlb_entry_ports_25_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_vpn_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_vpn_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_vpn_tlb_entry_ports_26_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_vpn_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_vpn_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_vpn_tlb_entry_ports_27_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_vpn_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_vpn_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_vpn_tlb_entry_ports_28_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_vpn_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_vpn_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_vpn_tlb_entry_ports_29_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_vpn_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_vpn_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_vpn_tlb_entry_ports_30_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_vpn_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_vpn_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_vpn_tlb_entry_ports_31_w_data = io_wport_bits_entry_vpn;
  assign tlb_entries_vpn_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_vpn_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_vpn_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_g__T_5_addr = 5'h0;
  assign tlb_entries_g__T_5_data = tlb_entries_g[tlb_entries_g__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_6_addr = 5'h1;
  assign tlb_entries_g__T_6_data = tlb_entries_g[tlb_entries_g__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_7_addr = 5'h2;
  assign tlb_entries_g__T_7_data = tlb_entries_g[tlb_entries_g__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_8_addr = 5'h3;
  assign tlb_entries_g__T_8_data = tlb_entries_g[tlb_entries_g__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_9_addr = 5'h4;
  assign tlb_entries_g__T_9_data = tlb_entries_g[tlb_entries_g__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_10_addr = 5'h5;
  assign tlb_entries_g__T_10_data = tlb_entries_g[tlb_entries_g__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_11_addr = 5'h6;
  assign tlb_entries_g__T_11_data = tlb_entries_g[tlb_entries_g__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_12_addr = 5'h7;
  assign tlb_entries_g__T_12_data = tlb_entries_g[tlb_entries_g__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_13_addr = 5'h8;
  assign tlb_entries_g__T_13_data = tlb_entries_g[tlb_entries_g__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_14_addr = 5'h9;
  assign tlb_entries_g__T_14_data = tlb_entries_g[tlb_entries_g__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_15_addr = 5'ha;
  assign tlb_entries_g__T_15_data = tlb_entries_g[tlb_entries_g__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_16_addr = 5'hb;
  assign tlb_entries_g__T_16_data = tlb_entries_g[tlb_entries_g__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_17_addr = 5'hc;
  assign tlb_entries_g__T_17_data = tlb_entries_g[tlb_entries_g__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_18_addr = 5'hd;
  assign tlb_entries_g__T_18_data = tlb_entries_g[tlb_entries_g__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_19_addr = 5'he;
  assign tlb_entries_g__T_19_data = tlb_entries_g[tlb_entries_g__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_20_addr = 5'hf;
  assign tlb_entries_g__T_20_data = tlb_entries_g[tlb_entries_g__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_21_addr = 5'h10;
  assign tlb_entries_g__T_21_data = tlb_entries_g[tlb_entries_g__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_22_addr = 5'h11;
  assign tlb_entries_g__T_22_data = tlb_entries_g[tlb_entries_g__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_23_addr = 5'h12;
  assign tlb_entries_g__T_23_data = tlb_entries_g[tlb_entries_g__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_24_addr = 5'h13;
  assign tlb_entries_g__T_24_data = tlb_entries_g[tlb_entries_g__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_25_addr = 5'h14;
  assign tlb_entries_g__T_25_data = tlb_entries_g[tlb_entries_g__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_26_addr = 5'h15;
  assign tlb_entries_g__T_26_data = tlb_entries_g[tlb_entries_g__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_27_addr = 5'h16;
  assign tlb_entries_g__T_27_data = tlb_entries_g[tlb_entries_g__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_28_addr = 5'h17;
  assign tlb_entries_g__T_28_data = tlb_entries_g[tlb_entries_g__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_29_addr = 5'h18;
  assign tlb_entries_g__T_29_data = tlb_entries_g[tlb_entries_g__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_30_addr = 5'h19;
  assign tlb_entries_g__T_30_data = tlb_entries_g[tlb_entries_g__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_31_addr = 5'h1a;
  assign tlb_entries_g__T_31_data = tlb_entries_g[tlb_entries_g__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_32_addr = 5'h1b;
  assign tlb_entries_g__T_32_data = tlb_entries_g[tlb_entries_g__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_33_addr = 5'h1c;
  assign tlb_entries_g__T_33_data = tlb_entries_g[tlb_entries_g__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_34_addr = 5'h1d;
  assign tlb_entries_g__T_34_data = tlb_entries_g[tlb_entries_g__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_35_addr = 5'h1e;
  assign tlb_entries_g__T_35_data = tlb_entries_g[tlb_entries_g__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_36_addr = 5'h1f;
  assign tlb_entries_g__T_36_data = tlb_entries_g[tlb_entries_g__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1546_addr = 5'h0;
  assign tlb_entries_g__T_1546_data = tlb_entries_g[tlb_entries_g__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1547_addr = 5'h1;
  assign tlb_entries_g__T_1547_data = tlb_entries_g[tlb_entries_g__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1548_addr = 5'h2;
  assign tlb_entries_g__T_1548_data = tlb_entries_g[tlb_entries_g__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1549_addr = 5'h3;
  assign tlb_entries_g__T_1549_data = tlb_entries_g[tlb_entries_g__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1550_addr = 5'h4;
  assign tlb_entries_g__T_1550_data = tlb_entries_g[tlb_entries_g__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1551_addr = 5'h5;
  assign tlb_entries_g__T_1551_data = tlb_entries_g[tlb_entries_g__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1552_addr = 5'h6;
  assign tlb_entries_g__T_1552_data = tlb_entries_g[tlb_entries_g__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1553_addr = 5'h7;
  assign tlb_entries_g__T_1553_data = tlb_entries_g[tlb_entries_g__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1554_addr = 5'h8;
  assign tlb_entries_g__T_1554_data = tlb_entries_g[tlb_entries_g__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1555_addr = 5'h9;
  assign tlb_entries_g__T_1555_data = tlb_entries_g[tlb_entries_g__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1556_addr = 5'ha;
  assign tlb_entries_g__T_1556_data = tlb_entries_g[tlb_entries_g__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1557_addr = 5'hb;
  assign tlb_entries_g__T_1557_data = tlb_entries_g[tlb_entries_g__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1558_addr = 5'hc;
  assign tlb_entries_g__T_1558_data = tlb_entries_g[tlb_entries_g__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1559_addr = 5'hd;
  assign tlb_entries_g__T_1559_data = tlb_entries_g[tlb_entries_g__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1560_addr = 5'he;
  assign tlb_entries_g__T_1560_data = tlb_entries_g[tlb_entries_g__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1561_addr = 5'hf;
  assign tlb_entries_g__T_1561_data = tlb_entries_g[tlb_entries_g__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1562_addr = 5'h10;
  assign tlb_entries_g__T_1562_data = tlb_entries_g[tlb_entries_g__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1563_addr = 5'h11;
  assign tlb_entries_g__T_1563_data = tlb_entries_g[tlb_entries_g__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1564_addr = 5'h12;
  assign tlb_entries_g__T_1564_data = tlb_entries_g[tlb_entries_g__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1565_addr = 5'h13;
  assign tlb_entries_g__T_1565_data = tlb_entries_g[tlb_entries_g__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1566_addr = 5'h14;
  assign tlb_entries_g__T_1566_data = tlb_entries_g[tlb_entries_g__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1567_addr = 5'h15;
  assign tlb_entries_g__T_1567_data = tlb_entries_g[tlb_entries_g__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1568_addr = 5'h16;
  assign tlb_entries_g__T_1568_data = tlb_entries_g[tlb_entries_g__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1569_addr = 5'h17;
  assign tlb_entries_g__T_1569_data = tlb_entries_g[tlb_entries_g__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1570_addr = 5'h18;
  assign tlb_entries_g__T_1570_data = tlb_entries_g[tlb_entries_g__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1571_addr = 5'h19;
  assign tlb_entries_g__T_1571_data = tlb_entries_g[tlb_entries_g__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1572_addr = 5'h1a;
  assign tlb_entries_g__T_1572_data = tlb_entries_g[tlb_entries_g__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1573_addr = 5'h1b;
  assign tlb_entries_g__T_1573_data = tlb_entries_g[tlb_entries_g__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1574_addr = 5'h1c;
  assign tlb_entries_g__T_1574_data = tlb_entries_g[tlb_entries_g__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1575_addr = 5'h1d;
  assign tlb_entries_g__T_1575_data = tlb_entries_g[tlb_entries_g__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1576_addr = 5'h1e;
  assign tlb_entries_g__T_1576_data = tlb_entries_g[tlb_entries_g__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g__T_1577_addr = 5'h1f;
  assign tlb_entries_g__T_1577_data = tlb_entries_g[tlb_entries_g__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_g_tlb_entry_ports_0_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_g_tlb_entry_ports_1_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_g_tlb_entry_ports_2_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_g_tlb_entry_ports_3_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_g_tlb_entry_ports_4_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_g_tlb_entry_ports_5_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_g_tlb_entry_ports_6_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_g_tlb_entry_ports_7_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_g_tlb_entry_ports_8_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_g_tlb_entry_ports_9_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_g_tlb_entry_ports_10_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_g_tlb_entry_ports_11_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_g_tlb_entry_ports_12_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_g_tlb_entry_ports_13_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_g_tlb_entry_ports_14_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_g_tlb_entry_ports_15_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_g_tlb_entry_ports_16_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_g_tlb_entry_ports_17_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_g_tlb_entry_ports_18_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_g_tlb_entry_ports_19_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_g_tlb_entry_ports_20_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_g_tlb_entry_ports_21_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_g_tlb_entry_ports_22_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_g_tlb_entry_ports_23_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_g_tlb_entry_ports_24_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_g_tlb_entry_ports_25_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_g_tlb_entry_ports_26_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_g_tlb_entry_ports_27_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_g_tlb_entry_ports_28_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_g_tlb_entry_ports_29_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_g_tlb_entry_ports_30_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_g_tlb_entry_ports_31_r_data = tlb_entries_g[tlb_entries_g_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_g_tlb_entry_ports_0_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_g_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_g_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_g_tlb_entry_ports_1_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_g_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_g_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_g_tlb_entry_ports_2_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_g_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_g_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_g_tlb_entry_ports_3_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_g_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_g_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_g_tlb_entry_ports_4_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_g_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_g_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_g_tlb_entry_ports_5_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_g_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_g_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_g_tlb_entry_ports_6_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_g_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_g_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_g_tlb_entry_ports_7_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_g_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_g_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_g_tlb_entry_ports_8_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_g_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_g_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_g_tlb_entry_ports_9_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_g_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_g_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_g_tlb_entry_ports_10_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_g_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_g_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_g_tlb_entry_ports_11_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_g_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_g_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_g_tlb_entry_ports_12_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_g_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_g_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_g_tlb_entry_ports_13_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_g_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_g_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_g_tlb_entry_ports_14_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_g_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_g_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_g_tlb_entry_ports_15_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_g_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_g_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_g_tlb_entry_ports_16_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_g_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_g_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_g_tlb_entry_ports_17_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_g_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_g_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_g_tlb_entry_ports_18_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_g_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_g_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_g_tlb_entry_ports_19_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_g_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_g_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_g_tlb_entry_ports_20_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_g_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_g_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_g_tlb_entry_ports_21_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_g_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_g_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_g_tlb_entry_ports_22_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_g_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_g_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_g_tlb_entry_ports_23_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_g_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_g_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_g_tlb_entry_ports_24_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_g_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_g_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_g_tlb_entry_ports_25_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_g_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_g_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_g_tlb_entry_ports_26_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_g_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_g_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_g_tlb_entry_ports_27_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_g_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_g_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_g_tlb_entry_ports_28_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_g_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_g_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_g_tlb_entry_ports_29_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_g_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_g_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_g_tlb_entry_ports_30_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_g_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_g_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_g_tlb_entry_ports_31_w_data = io_wport_bits_entry_g;
  assign tlb_entries_g_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_g_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_g_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_asid__T_5_addr = 5'h0;
  assign tlb_entries_asid__T_5_data = tlb_entries_asid[tlb_entries_asid__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_6_addr = 5'h1;
  assign tlb_entries_asid__T_6_data = tlb_entries_asid[tlb_entries_asid__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_7_addr = 5'h2;
  assign tlb_entries_asid__T_7_data = tlb_entries_asid[tlb_entries_asid__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_8_addr = 5'h3;
  assign tlb_entries_asid__T_8_data = tlb_entries_asid[tlb_entries_asid__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_9_addr = 5'h4;
  assign tlb_entries_asid__T_9_data = tlb_entries_asid[tlb_entries_asid__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_10_addr = 5'h5;
  assign tlb_entries_asid__T_10_data = tlb_entries_asid[tlb_entries_asid__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_11_addr = 5'h6;
  assign tlb_entries_asid__T_11_data = tlb_entries_asid[tlb_entries_asid__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_12_addr = 5'h7;
  assign tlb_entries_asid__T_12_data = tlb_entries_asid[tlb_entries_asid__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_13_addr = 5'h8;
  assign tlb_entries_asid__T_13_data = tlb_entries_asid[tlb_entries_asid__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_14_addr = 5'h9;
  assign tlb_entries_asid__T_14_data = tlb_entries_asid[tlb_entries_asid__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_15_addr = 5'ha;
  assign tlb_entries_asid__T_15_data = tlb_entries_asid[tlb_entries_asid__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_16_addr = 5'hb;
  assign tlb_entries_asid__T_16_data = tlb_entries_asid[tlb_entries_asid__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_17_addr = 5'hc;
  assign tlb_entries_asid__T_17_data = tlb_entries_asid[tlb_entries_asid__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_18_addr = 5'hd;
  assign tlb_entries_asid__T_18_data = tlb_entries_asid[tlb_entries_asid__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_19_addr = 5'he;
  assign tlb_entries_asid__T_19_data = tlb_entries_asid[tlb_entries_asid__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_20_addr = 5'hf;
  assign tlb_entries_asid__T_20_data = tlb_entries_asid[tlb_entries_asid__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_21_addr = 5'h10;
  assign tlb_entries_asid__T_21_data = tlb_entries_asid[tlb_entries_asid__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_22_addr = 5'h11;
  assign tlb_entries_asid__T_22_data = tlb_entries_asid[tlb_entries_asid__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_23_addr = 5'h12;
  assign tlb_entries_asid__T_23_data = tlb_entries_asid[tlb_entries_asid__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_24_addr = 5'h13;
  assign tlb_entries_asid__T_24_data = tlb_entries_asid[tlb_entries_asid__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_25_addr = 5'h14;
  assign tlb_entries_asid__T_25_data = tlb_entries_asid[tlb_entries_asid__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_26_addr = 5'h15;
  assign tlb_entries_asid__T_26_data = tlb_entries_asid[tlb_entries_asid__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_27_addr = 5'h16;
  assign tlb_entries_asid__T_27_data = tlb_entries_asid[tlb_entries_asid__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_28_addr = 5'h17;
  assign tlb_entries_asid__T_28_data = tlb_entries_asid[tlb_entries_asid__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_29_addr = 5'h18;
  assign tlb_entries_asid__T_29_data = tlb_entries_asid[tlb_entries_asid__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_30_addr = 5'h19;
  assign tlb_entries_asid__T_30_data = tlb_entries_asid[tlb_entries_asid__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_31_addr = 5'h1a;
  assign tlb_entries_asid__T_31_data = tlb_entries_asid[tlb_entries_asid__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_32_addr = 5'h1b;
  assign tlb_entries_asid__T_32_data = tlb_entries_asid[tlb_entries_asid__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_33_addr = 5'h1c;
  assign tlb_entries_asid__T_33_data = tlb_entries_asid[tlb_entries_asid__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_34_addr = 5'h1d;
  assign tlb_entries_asid__T_34_data = tlb_entries_asid[tlb_entries_asid__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_35_addr = 5'h1e;
  assign tlb_entries_asid__T_35_data = tlb_entries_asid[tlb_entries_asid__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_36_addr = 5'h1f;
  assign tlb_entries_asid__T_36_data = tlb_entries_asid[tlb_entries_asid__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1546_addr = 5'h0;
  assign tlb_entries_asid__T_1546_data = tlb_entries_asid[tlb_entries_asid__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1547_addr = 5'h1;
  assign tlb_entries_asid__T_1547_data = tlb_entries_asid[tlb_entries_asid__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1548_addr = 5'h2;
  assign tlb_entries_asid__T_1548_data = tlb_entries_asid[tlb_entries_asid__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1549_addr = 5'h3;
  assign tlb_entries_asid__T_1549_data = tlb_entries_asid[tlb_entries_asid__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1550_addr = 5'h4;
  assign tlb_entries_asid__T_1550_data = tlb_entries_asid[tlb_entries_asid__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1551_addr = 5'h5;
  assign tlb_entries_asid__T_1551_data = tlb_entries_asid[tlb_entries_asid__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1552_addr = 5'h6;
  assign tlb_entries_asid__T_1552_data = tlb_entries_asid[tlb_entries_asid__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1553_addr = 5'h7;
  assign tlb_entries_asid__T_1553_data = tlb_entries_asid[tlb_entries_asid__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1554_addr = 5'h8;
  assign tlb_entries_asid__T_1554_data = tlb_entries_asid[tlb_entries_asid__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1555_addr = 5'h9;
  assign tlb_entries_asid__T_1555_data = tlb_entries_asid[tlb_entries_asid__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1556_addr = 5'ha;
  assign tlb_entries_asid__T_1556_data = tlb_entries_asid[tlb_entries_asid__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1557_addr = 5'hb;
  assign tlb_entries_asid__T_1557_data = tlb_entries_asid[tlb_entries_asid__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1558_addr = 5'hc;
  assign tlb_entries_asid__T_1558_data = tlb_entries_asid[tlb_entries_asid__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1559_addr = 5'hd;
  assign tlb_entries_asid__T_1559_data = tlb_entries_asid[tlb_entries_asid__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1560_addr = 5'he;
  assign tlb_entries_asid__T_1560_data = tlb_entries_asid[tlb_entries_asid__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1561_addr = 5'hf;
  assign tlb_entries_asid__T_1561_data = tlb_entries_asid[tlb_entries_asid__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1562_addr = 5'h10;
  assign tlb_entries_asid__T_1562_data = tlb_entries_asid[tlb_entries_asid__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1563_addr = 5'h11;
  assign tlb_entries_asid__T_1563_data = tlb_entries_asid[tlb_entries_asid__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1564_addr = 5'h12;
  assign tlb_entries_asid__T_1564_data = tlb_entries_asid[tlb_entries_asid__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1565_addr = 5'h13;
  assign tlb_entries_asid__T_1565_data = tlb_entries_asid[tlb_entries_asid__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1566_addr = 5'h14;
  assign tlb_entries_asid__T_1566_data = tlb_entries_asid[tlb_entries_asid__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1567_addr = 5'h15;
  assign tlb_entries_asid__T_1567_data = tlb_entries_asid[tlb_entries_asid__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1568_addr = 5'h16;
  assign tlb_entries_asid__T_1568_data = tlb_entries_asid[tlb_entries_asid__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1569_addr = 5'h17;
  assign tlb_entries_asid__T_1569_data = tlb_entries_asid[tlb_entries_asid__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1570_addr = 5'h18;
  assign tlb_entries_asid__T_1570_data = tlb_entries_asid[tlb_entries_asid__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1571_addr = 5'h19;
  assign tlb_entries_asid__T_1571_data = tlb_entries_asid[tlb_entries_asid__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1572_addr = 5'h1a;
  assign tlb_entries_asid__T_1572_data = tlb_entries_asid[tlb_entries_asid__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1573_addr = 5'h1b;
  assign tlb_entries_asid__T_1573_data = tlb_entries_asid[tlb_entries_asid__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1574_addr = 5'h1c;
  assign tlb_entries_asid__T_1574_data = tlb_entries_asid[tlb_entries_asid__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1575_addr = 5'h1d;
  assign tlb_entries_asid__T_1575_data = tlb_entries_asid[tlb_entries_asid__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1576_addr = 5'h1e;
  assign tlb_entries_asid__T_1576_data = tlb_entries_asid[tlb_entries_asid__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid__T_1577_addr = 5'h1f;
  assign tlb_entries_asid__T_1577_data = tlb_entries_asid[tlb_entries_asid__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_asid_tlb_entry_ports_0_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_asid_tlb_entry_ports_1_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_asid_tlb_entry_ports_2_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_asid_tlb_entry_ports_3_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_asid_tlb_entry_ports_4_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_asid_tlb_entry_ports_5_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_asid_tlb_entry_ports_6_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_asid_tlb_entry_ports_7_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_asid_tlb_entry_ports_8_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_asid_tlb_entry_ports_9_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_asid_tlb_entry_ports_10_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_asid_tlb_entry_ports_11_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_asid_tlb_entry_ports_12_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_asid_tlb_entry_ports_13_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_asid_tlb_entry_ports_14_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_asid_tlb_entry_ports_15_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_asid_tlb_entry_ports_16_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_asid_tlb_entry_ports_17_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_asid_tlb_entry_ports_18_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_asid_tlb_entry_ports_19_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_asid_tlb_entry_ports_20_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_asid_tlb_entry_ports_21_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_asid_tlb_entry_ports_22_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_asid_tlb_entry_ports_23_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_asid_tlb_entry_ports_24_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_asid_tlb_entry_ports_25_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_asid_tlb_entry_ports_26_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_asid_tlb_entry_ports_27_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_asid_tlb_entry_ports_28_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_asid_tlb_entry_ports_29_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_asid_tlb_entry_ports_30_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_asid_tlb_entry_ports_31_r_data = tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_asid_tlb_entry_ports_0_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_asid_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_asid_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_asid_tlb_entry_ports_1_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_asid_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_asid_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_asid_tlb_entry_ports_2_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_asid_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_asid_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_asid_tlb_entry_ports_3_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_asid_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_asid_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_asid_tlb_entry_ports_4_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_asid_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_asid_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_asid_tlb_entry_ports_5_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_asid_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_asid_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_asid_tlb_entry_ports_6_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_asid_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_asid_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_asid_tlb_entry_ports_7_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_asid_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_asid_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_asid_tlb_entry_ports_8_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_asid_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_asid_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_asid_tlb_entry_ports_9_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_asid_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_asid_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_asid_tlb_entry_ports_10_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_asid_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_asid_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_asid_tlb_entry_ports_11_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_asid_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_asid_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_asid_tlb_entry_ports_12_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_asid_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_asid_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_asid_tlb_entry_ports_13_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_asid_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_asid_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_asid_tlb_entry_ports_14_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_asid_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_asid_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_asid_tlb_entry_ports_15_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_asid_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_asid_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_asid_tlb_entry_ports_16_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_asid_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_asid_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_asid_tlb_entry_ports_17_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_asid_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_asid_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_asid_tlb_entry_ports_18_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_asid_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_asid_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_asid_tlb_entry_ports_19_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_asid_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_asid_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_asid_tlb_entry_ports_20_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_asid_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_asid_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_asid_tlb_entry_ports_21_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_asid_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_asid_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_asid_tlb_entry_ports_22_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_asid_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_asid_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_asid_tlb_entry_ports_23_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_asid_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_asid_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_asid_tlb_entry_ports_24_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_asid_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_asid_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_asid_tlb_entry_ports_25_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_asid_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_asid_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_asid_tlb_entry_ports_26_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_asid_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_asid_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_asid_tlb_entry_ports_27_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_asid_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_asid_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_asid_tlb_entry_ports_28_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_asid_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_asid_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_asid_tlb_entry_ports_29_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_asid_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_asid_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_asid_tlb_entry_ports_30_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_asid_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_asid_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_asid_tlb_entry_ports_31_w_data = io_wport_bits_entry_asid;
  assign tlb_entries_asid_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_asid_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_asid_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p0_pfn__T_5_addr = 5'h0;
  assign tlb_entries_p0_pfn__T_5_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_6_addr = 5'h1;
  assign tlb_entries_p0_pfn__T_6_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_7_addr = 5'h2;
  assign tlb_entries_p0_pfn__T_7_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_8_addr = 5'h3;
  assign tlb_entries_p0_pfn__T_8_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_9_addr = 5'h4;
  assign tlb_entries_p0_pfn__T_9_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_10_addr = 5'h5;
  assign tlb_entries_p0_pfn__T_10_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_11_addr = 5'h6;
  assign tlb_entries_p0_pfn__T_11_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_12_addr = 5'h7;
  assign tlb_entries_p0_pfn__T_12_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_13_addr = 5'h8;
  assign tlb_entries_p0_pfn__T_13_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_14_addr = 5'h9;
  assign tlb_entries_p0_pfn__T_14_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_15_addr = 5'ha;
  assign tlb_entries_p0_pfn__T_15_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_16_addr = 5'hb;
  assign tlb_entries_p0_pfn__T_16_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_17_addr = 5'hc;
  assign tlb_entries_p0_pfn__T_17_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_18_addr = 5'hd;
  assign tlb_entries_p0_pfn__T_18_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_19_addr = 5'he;
  assign tlb_entries_p0_pfn__T_19_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_20_addr = 5'hf;
  assign tlb_entries_p0_pfn__T_20_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_21_addr = 5'h10;
  assign tlb_entries_p0_pfn__T_21_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_22_addr = 5'h11;
  assign tlb_entries_p0_pfn__T_22_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_23_addr = 5'h12;
  assign tlb_entries_p0_pfn__T_23_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_24_addr = 5'h13;
  assign tlb_entries_p0_pfn__T_24_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_25_addr = 5'h14;
  assign tlb_entries_p0_pfn__T_25_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_26_addr = 5'h15;
  assign tlb_entries_p0_pfn__T_26_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_27_addr = 5'h16;
  assign tlb_entries_p0_pfn__T_27_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_28_addr = 5'h17;
  assign tlb_entries_p0_pfn__T_28_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_29_addr = 5'h18;
  assign tlb_entries_p0_pfn__T_29_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_30_addr = 5'h19;
  assign tlb_entries_p0_pfn__T_30_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_31_addr = 5'h1a;
  assign tlb_entries_p0_pfn__T_31_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_32_addr = 5'h1b;
  assign tlb_entries_p0_pfn__T_32_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_33_addr = 5'h1c;
  assign tlb_entries_p0_pfn__T_33_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_34_addr = 5'h1d;
  assign tlb_entries_p0_pfn__T_34_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_35_addr = 5'h1e;
  assign tlb_entries_p0_pfn__T_35_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_36_addr = 5'h1f;
  assign tlb_entries_p0_pfn__T_36_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1546_addr = 5'h0;
  assign tlb_entries_p0_pfn__T_1546_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1547_addr = 5'h1;
  assign tlb_entries_p0_pfn__T_1547_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1548_addr = 5'h2;
  assign tlb_entries_p0_pfn__T_1548_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1549_addr = 5'h3;
  assign tlb_entries_p0_pfn__T_1549_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1550_addr = 5'h4;
  assign tlb_entries_p0_pfn__T_1550_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1551_addr = 5'h5;
  assign tlb_entries_p0_pfn__T_1551_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1552_addr = 5'h6;
  assign tlb_entries_p0_pfn__T_1552_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1553_addr = 5'h7;
  assign tlb_entries_p0_pfn__T_1553_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1554_addr = 5'h8;
  assign tlb_entries_p0_pfn__T_1554_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1555_addr = 5'h9;
  assign tlb_entries_p0_pfn__T_1555_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1556_addr = 5'ha;
  assign tlb_entries_p0_pfn__T_1556_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1557_addr = 5'hb;
  assign tlb_entries_p0_pfn__T_1557_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1558_addr = 5'hc;
  assign tlb_entries_p0_pfn__T_1558_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1559_addr = 5'hd;
  assign tlb_entries_p0_pfn__T_1559_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1560_addr = 5'he;
  assign tlb_entries_p0_pfn__T_1560_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1561_addr = 5'hf;
  assign tlb_entries_p0_pfn__T_1561_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1562_addr = 5'h10;
  assign tlb_entries_p0_pfn__T_1562_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1563_addr = 5'h11;
  assign tlb_entries_p0_pfn__T_1563_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1564_addr = 5'h12;
  assign tlb_entries_p0_pfn__T_1564_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1565_addr = 5'h13;
  assign tlb_entries_p0_pfn__T_1565_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1566_addr = 5'h14;
  assign tlb_entries_p0_pfn__T_1566_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1567_addr = 5'h15;
  assign tlb_entries_p0_pfn__T_1567_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1568_addr = 5'h16;
  assign tlb_entries_p0_pfn__T_1568_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1569_addr = 5'h17;
  assign tlb_entries_p0_pfn__T_1569_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1570_addr = 5'h18;
  assign tlb_entries_p0_pfn__T_1570_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1571_addr = 5'h19;
  assign tlb_entries_p0_pfn__T_1571_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1572_addr = 5'h1a;
  assign tlb_entries_p0_pfn__T_1572_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1573_addr = 5'h1b;
  assign tlb_entries_p0_pfn__T_1573_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1574_addr = 5'h1c;
  assign tlb_entries_p0_pfn__T_1574_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1575_addr = 5'h1d;
  assign tlb_entries_p0_pfn__T_1575_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1576_addr = 5'h1e;
  assign tlb_entries_p0_pfn__T_1576_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn__T_1577_addr = 5'h1f;
  assign tlb_entries_p0_pfn__T_1577_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p0_pfn_tlb_entry_ports_0_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p0_pfn_tlb_entry_ports_1_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p0_pfn_tlb_entry_ports_2_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p0_pfn_tlb_entry_ports_3_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p0_pfn_tlb_entry_ports_4_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p0_pfn_tlb_entry_ports_5_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p0_pfn_tlb_entry_ports_6_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p0_pfn_tlb_entry_ports_7_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p0_pfn_tlb_entry_ports_8_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p0_pfn_tlb_entry_ports_9_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p0_pfn_tlb_entry_ports_10_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p0_pfn_tlb_entry_ports_11_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p0_pfn_tlb_entry_ports_12_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p0_pfn_tlb_entry_ports_13_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p0_pfn_tlb_entry_ports_14_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p0_pfn_tlb_entry_ports_15_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p0_pfn_tlb_entry_ports_16_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p0_pfn_tlb_entry_ports_17_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p0_pfn_tlb_entry_ports_18_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p0_pfn_tlb_entry_ports_19_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p0_pfn_tlb_entry_ports_20_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p0_pfn_tlb_entry_ports_21_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p0_pfn_tlb_entry_ports_22_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p0_pfn_tlb_entry_ports_23_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p0_pfn_tlb_entry_ports_24_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p0_pfn_tlb_entry_ports_25_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p0_pfn_tlb_entry_ports_26_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p0_pfn_tlb_entry_ports_27_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p0_pfn_tlb_entry_ports_28_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p0_pfn_tlb_entry_ports_29_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p0_pfn_tlb_entry_ports_30_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p0_pfn_tlb_entry_ports_31_r_data = tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_pfn_tlb_entry_ports_0_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p0_pfn_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p0_pfn_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p0_pfn_tlb_entry_ports_1_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p0_pfn_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p0_pfn_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p0_pfn_tlb_entry_ports_2_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p0_pfn_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p0_pfn_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p0_pfn_tlb_entry_ports_3_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p0_pfn_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p0_pfn_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p0_pfn_tlb_entry_ports_4_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p0_pfn_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p0_pfn_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p0_pfn_tlb_entry_ports_5_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p0_pfn_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p0_pfn_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p0_pfn_tlb_entry_ports_6_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p0_pfn_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p0_pfn_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p0_pfn_tlb_entry_ports_7_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p0_pfn_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p0_pfn_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p0_pfn_tlb_entry_ports_8_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p0_pfn_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p0_pfn_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p0_pfn_tlb_entry_ports_9_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p0_pfn_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p0_pfn_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p0_pfn_tlb_entry_ports_10_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p0_pfn_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p0_pfn_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p0_pfn_tlb_entry_ports_11_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p0_pfn_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p0_pfn_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p0_pfn_tlb_entry_ports_12_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p0_pfn_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p0_pfn_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p0_pfn_tlb_entry_ports_13_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p0_pfn_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p0_pfn_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p0_pfn_tlb_entry_ports_14_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p0_pfn_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p0_pfn_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p0_pfn_tlb_entry_ports_15_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p0_pfn_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p0_pfn_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p0_pfn_tlb_entry_ports_16_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p0_pfn_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p0_pfn_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p0_pfn_tlb_entry_ports_17_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p0_pfn_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p0_pfn_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p0_pfn_tlb_entry_ports_18_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p0_pfn_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p0_pfn_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p0_pfn_tlb_entry_ports_19_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p0_pfn_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p0_pfn_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p0_pfn_tlb_entry_ports_20_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p0_pfn_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p0_pfn_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p0_pfn_tlb_entry_ports_21_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p0_pfn_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p0_pfn_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p0_pfn_tlb_entry_ports_22_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p0_pfn_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p0_pfn_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p0_pfn_tlb_entry_ports_23_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p0_pfn_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p0_pfn_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p0_pfn_tlb_entry_ports_24_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p0_pfn_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p0_pfn_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p0_pfn_tlb_entry_ports_25_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p0_pfn_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p0_pfn_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p0_pfn_tlb_entry_ports_26_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p0_pfn_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p0_pfn_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p0_pfn_tlb_entry_ports_27_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p0_pfn_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p0_pfn_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p0_pfn_tlb_entry_ports_28_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p0_pfn_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p0_pfn_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p0_pfn_tlb_entry_ports_29_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p0_pfn_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p0_pfn_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p0_pfn_tlb_entry_ports_30_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p0_pfn_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p0_pfn_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p0_pfn_tlb_entry_ports_31_w_data = io_wport_bits_entry_p0_pfn;
  assign tlb_entries_p0_pfn_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p0_pfn_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p0_pfn_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p0_c__T_5_addr = 5'h0;
  assign tlb_entries_p0_c__T_5_data = tlb_entries_p0_c[tlb_entries_p0_c__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_6_addr = 5'h1;
  assign tlb_entries_p0_c__T_6_data = tlb_entries_p0_c[tlb_entries_p0_c__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_7_addr = 5'h2;
  assign tlb_entries_p0_c__T_7_data = tlb_entries_p0_c[tlb_entries_p0_c__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_8_addr = 5'h3;
  assign tlb_entries_p0_c__T_8_data = tlb_entries_p0_c[tlb_entries_p0_c__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_9_addr = 5'h4;
  assign tlb_entries_p0_c__T_9_data = tlb_entries_p0_c[tlb_entries_p0_c__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_10_addr = 5'h5;
  assign tlb_entries_p0_c__T_10_data = tlb_entries_p0_c[tlb_entries_p0_c__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_11_addr = 5'h6;
  assign tlb_entries_p0_c__T_11_data = tlb_entries_p0_c[tlb_entries_p0_c__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_12_addr = 5'h7;
  assign tlb_entries_p0_c__T_12_data = tlb_entries_p0_c[tlb_entries_p0_c__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_13_addr = 5'h8;
  assign tlb_entries_p0_c__T_13_data = tlb_entries_p0_c[tlb_entries_p0_c__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_14_addr = 5'h9;
  assign tlb_entries_p0_c__T_14_data = tlb_entries_p0_c[tlb_entries_p0_c__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_15_addr = 5'ha;
  assign tlb_entries_p0_c__T_15_data = tlb_entries_p0_c[tlb_entries_p0_c__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_16_addr = 5'hb;
  assign tlb_entries_p0_c__T_16_data = tlb_entries_p0_c[tlb_entries_p0_c__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_17_addr = 5'hc;
  assign tlb_entries_p0_c__T_17_data = tlb_entries_p0_c[tlb_entries_p0_c__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_18_addr = 5'hd;
  assign tlb_entries_p0_c__T_18_data = tlb_entries_p0_c[tlb_entries_p0_c__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_19_addr = 5'he;
  assign tlb_entries_p0_c__T_19_data = tlb_entries_p0_c[tlb_entries_p0_c__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_20_addr = 5'hf;
  assign tlb_entries_p0_c__T_20_data = tlb_entries_p0_c[tlb_entries_p0_c__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_21_addr = 5'h10;
  assign tlb_entries_p0_c__T_21_data = tlb_entries_p0_c[tlb_entries_p0_c__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_22_addr = 5'h11;
  assign tlb_entries_p0_c__T_22_data = tlb_entries_p0_c[tlb_entries_p0_c__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_23_addr = 5'h12;
  assign tlb_entries_p0_c__T_23_data = tlb_entries_p0_c[tlb_entries_p0_c__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_24_addr = 5'h13;
  assign tlb_entries_p0_c__T_24_data = tlb_entries_p0_c[tlb_entries_p0_c__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_25_addr = 5'h14;
  assign tlb_entries_p0_c__T_25_data = tlb_entries_p0_c[tlb_entries_p0_c__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_26_addr = 5'h15;
  assign tlb_entries_p0_c__T_26_data = tlb_entries_p0_c[tlb_entries_p0_c__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_27_addr = 5'h16;
  assign tlb_entries_p0_c__T_27_data = tlb_entries_p0_c[tlb_entries_p0_c__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_28_addr = 5'h17;
  assign tlb_entries_p0_c__T_28_data = tlb_entries_p0_c[tlb_entries_p0_c__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_29_addr = 5'h18;
  assign tlb_entries_p0_c__T_29_data = tlb_entries_p0_c[tlb_entries_p0_c__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_30_addr = 5'h19;
  assign tlb_entries_p0_c__T_30_data = tlb_entries_p0_c[tlb_entries_p0_c__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_31_addr = 5'h1a;
  assign tlb_entries_p0_c__T_31_data = tlb_entries_p0_c[tlb_entries_p0_c__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_32_addr = 5'h1b;
  assign tlb_entries_p0_c__T_32_data = tlb_entries_p0_c[tlb_entries_p0_c__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_33_addr = 5'h1c;
  assign tlb_entries_p0_c__T_33_data = tlb_entries_p0_c[tlb_entries_p0_c__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_34_addr = 5'h1d;
  assign tlb_entries_p0_c__T_34_data = tlb_entries_p0_c[tlb_entries_p0_c__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_35_addr = 5'h1e;
  assign tlb_entries_p0_c__T_35_data = tlb_entries_p0_c[tlb_entries_p0_c__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_36_addr = 5'h1f;
  assign tlb_entries_p0_c__T_36_data = tlb_entries_p0_c[tlb_entries_p0_c__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1546_addr = 5'h0;
  assign tlb_entries_p0_c__T_1546_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1547_addr = 5'h1;
  assign tlb_entries_p0_c__T_1547_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1548_addr = 5'h2;
  assign tlb_entries_p0_c__T_1548_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1549_addr = 5'h3;
  assign tlb_entries_p0_c__T_1549_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1550_addr = 5'h4;
  assign tlb_entries_p0_c__T_1550_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1551_addr = 5'h5;
  assign tlb_entries_p0_c__T_1551_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1552_addr = 5'h6;
  assign tlb_entries_p0_c__T_1552_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1553_addr = 5'h7;
  assign tlb_entries_p0_c__T_1553_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1554_addr = 5'h8;
  assign tlb_entries_p0_c__T_1554_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1555_addr = 5'h9;
  assign tlb_entries_p0_c__T_1555_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1556_addr = 5'ha;
  assign tlb_entries_p0_c__T_1556_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1557_addr = 5'hb;
  assign tlb_entries_p0_c__T_1557_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1558_addr = 5'hc;
  assign tlb_entries_p0_c__T_1558_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1559_addr = 5'hd;
  assign tlb_entries_p0_c__T_1559_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1560_addr = 5'he;
  assign tlb_entries_p0_c__T_1560_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1561_addr = 5'hf;
  assign tlb_entries_p0_c__T_1561_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1562_addr = 5'h10;
  assign tlb_entries_p0_c__T_1562_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1563_addr = 5'h11;
  assign tlb_entries_p0_c__T_1563_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1564_addr = 5'h12;
  assign tlb_entries_p0_c__T_1564_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1565_addr = 5'h13;
  assign tlb_entries_p0_c__T_1565_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1566_addr = 5'h14;
  assign tlb_entries_p0_c__T_1566_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1567_addr = 5'h15;
  assign tlb_entries_p0_c__T_1567_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1568_addr = 5'h16;
  assign tlb_entries_p0_c__T_1568_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1569_addr = 5'h17;
  assign tlb_entries_p0_c__T_1569_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1570_addr = 5'h18;
  assign tlb_entries_p0_c__T_1570_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1571_addr = 5'h19;
  assign tlb_entries_p0_c__T_1571_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1572_addr = 5'h1a;
  assign tlb_entries_p0_c__T_1572_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1573_addr = 5'h1b;
  assign tlb_entries_p0_c__T_1573_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1574_addr = 5'h1c;
  assign tlb_entries_p0_c__T_1574_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1575_addr = 5'h1d;
  assign tlb_entries_p0_c__T_1575_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1576_addr = 5'h1e;
  assign tlb_entries_p0_c__T_1576_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c__T_1577_addr = 5'h1f;
  assign tlb_entries_p0_c__T_1577_data = tlb_entries_p0_c[tlb_entries_p0_c__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p0_c_tlb_entry_ports_0_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p0_c_tlb_entry_ports_1_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p0_c_tlb_entry_ports_2_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p0_c_tlb_entry_ports_3_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p0_c_tlb_entry_ports_4_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p0_c_tlb_entry_ports_5_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p0_c_tlb_entry_ports_6_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p0_c_tlb_entry_ports_7_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p0_c_tlb_entry_ports_8_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p0_c_tlb_entry_ports_9_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p0_c_tlb_entry_ports_10_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p0_c_tlb_entry_ports_11_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p0_c_tlb_entry_ports_12_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p0_c_tlb_entry_ports_13_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p0_c_tlb_entry_ports_14_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p0_c_tlb_entry_ports_15_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p0_c_tlb_entry_ports_16_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p0_c_tlb_entry_ports_17_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p0_c_tlb_entry_ports_18_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p0_c_tlb_entry_ports_19_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p0_c_tlb_entry_ports_20_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p0_c_tlb_entry_ports_21_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p0_c_tlb_entry_ports_22_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p0_c_tlb_entry_ports_23_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p0_c_tlb_entry_ports_24_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p0_c_tlb_entry_ports_25_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p0_c_tlb_entry_ports_26_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p0_c_tlb_entry_ports_27_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p0_c_tlb_entry_ports_28_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p0_c_tlb_entry_ports_29_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p0_c_tlb_entry_ports_30_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p0_c_tlb_entry_ports_31_r_data = tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_c_tlb_entry_ports_0_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p0_c_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p0_c_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p0_c_tlb_entry_ports_1_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p0_c_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p0_c_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p0_c_tlb_entry_ports_2_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p0_c_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p0_c_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p0_c_tlb_entry_ports_3_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p0_c_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p0_c_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p0_c_tlb_entry_ports_4_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p0_c_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p0_c_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p0_c_tlb_entry_ports_5_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p0_c_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p0_c_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p0_c_tlb_entry_ports_6_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p0_c_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p0_c_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p0_c_tlb_entry_ports_7_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p0_c_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p0_c_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p0_c_tlb_entry_ports_8_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p0_c_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p0_c_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p0_c_tlb_entry_ports_9_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p0_c_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p0_c_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p0_c_tlb_entry_ports_10_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p0_c_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p0_c_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p0_c_tlb_entry_ports_11_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p0_c_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p0_c_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p0_c_tlb_entry_ports_12_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p0_c_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p0_c_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p0_c_tlb_entry_ports_13_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p0_c_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p0_c_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p0_c_tlb_entry_ports_14_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p0_c_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p0_c_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p0_c_tlb_entry_ports_15_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p0_c_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p0_c_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p0_c_tlb_entry_ports_16_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p0_c_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p0_c_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p0_c_tlb_entry_ports_17_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p0_c_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p0_c_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p0_c_tlb_entry_ports_18_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p0_c_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p0_c_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p0_c_tlb_entry_ports_19_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p0_c_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p0_c_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p0_c_tlb_entry_ports_20_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p0_c_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p0_c_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p0_c_tlb_entry_ports_21_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p0_c_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p0_c_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p0_c_tlb_entry_ports_22_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p0_c_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p0_c_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p0_c_tlb_entry_ports_23_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p0_c_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p0_c_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p0_c_tlb_entry_ports_24_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p0_c_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p0_c_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p0_c_tlb_entry_ports_25_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p0_c_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p0_c_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p0_c_tlb_entry_ports_26_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p0_c_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p0_c_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p0_c_tlb_entry_ports_27_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p0_c_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p0_c_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p0_c_tlb_entry_ports_28_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p0_c_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p0_c_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p0_c_tlb_entry_ports_29_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p0_c_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p0_c_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p0_c_tlb_entry_ports_30_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p0_c_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p0_c_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p0_c_tlb_entry_ports_31_w_data = io_wport_bits_entry_p0_c;
  assign tlb_entries_p0_c_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p0_c_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p0_c_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p0_d__T_5_addr = 5'h0;
  assign tlb_entries_p0_d__T_5_data = tlb_entries_p0_d[tlb_entries_p0_d__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_6_addr = 5'h1;
  assign tlb_entries_p0_d__T_6_data = tlb_entries_p0_d[tlb_entries_p0_d__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_7_addr = 5'h2;
  assign tlb_entries_p0_d__T_7_data = tlb_entries_p0_d[tlb_entries_p0_d__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_8_addr = 5'h3;
  assign tlb_entries_p0_d__T_8_data = tlb_entries_p0_d[tlb_entries_p0_d__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_9_addr = 5'h4;
  assign tlb_entries_p0_d__T_9_data = tlb_entries_p0_d[tlb_entries_p0_d__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_10_addr = 5'h5;
  assign tlb_entries_p0_d__T_10_data = tlb_entries_p0_d[tlb_entries_p0_d__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_11_addr = 5'h6;
  assign tlb_entries_p0_d__T_11_data = tlb_entries_p0_d[tlb_entries_p0_d__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_12_addr = 5'h7;
  assign tlb_entries_p0_d__T_12_data = tlb_entries_p0_d[tlb_entries_p0_d__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_13_addr = 5'h8;
  assign tlb_entries_p0_d__T_13_data = tlb_entries_p0_d[tlb_entries_p0_d__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_14_addr = 5'h9;
  assign tlb_entries_p0_d__T_14_data = tlb_entries_p0_d[tlb_entries_p0_d__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_15_addr = 5'ha;
  assign tlb_entries_p0_d__T_15_data = tlb_entries_p0_d[tlb_entries_p0_d__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_16_addr = 5'hb;
  assign tlb_entries_p0_d__T_16_data = tlb_entries_p0_d[tlb_entries_p0_d__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_17_addr = 5'hc;
  assign tlb_entries_p0_d__T_17_data = tlb_entries_p0_d[tlb_entries_p0_d__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_18_addr = 5'hd;
  assign tlb_entries_p0_d__T_18_data = tlb_entries_p0_d[tlb_entries_p0_d__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_19_addr = 5'he;
  assign tlb_entries_p0_d__T_19_data = tlb_entries_p0_d[tlb_entries_p0_d__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_20_addr = 5'hf;
  assign tlb_entries_p0_d__T_20_data = tlb_entries_p0_d[tlb_entries_p0_d__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_21_addr = 5'h10;
  assign tlb_entries_p0_d__T_21_data = tlb_entries_p0_d[tlb_entries_p0_d__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_22_addr = 5'h11;
  assign tlb_entries_p0_d__T_22_data = tlb_entries_p0_d[tlb_entries_p0_d__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_23_addr = 5'h12;
  assign tlb_entries_p0_d__T_23_data = tlb_entries_p0_d[tlb_entries_p0_d__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_24_addr = 5'h13;
  assign tlb_entries_p0_d__T_24_data = tlb_entries_p0_d[tlb_entries_p0_d__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_25_addr = 5'h14;
  assign tlb_entries_p0_d__T_25_data = tlb_entries_p0_d[tlb_entries_p0_d__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_26_addr = 5'h15;
  assign tlb_entries_p0_d__T_26_data = tlb_entries_p0_d[tlb_entries_p0_d__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_27_addr = 5'h16;
  assign tlb_entries_p0_d__T_27_data = tlb_entries_p0_d[tlb_entries_p0_d__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_28_addr = 5'h17;
  assign tlb_entries_p0_d__T_28_data = tlb_entries_p0_d[tlb_entries_p0_d__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_29_addr = 5'h18;
  assign tlb_entries_p0_d__T_29_data = tlb_entries_p0_d[tlb_entries_p0_d__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_30_addr = 5'h19;
  assign tlb_entries_p0_d__T_30_data = tlb_entries_p0_d[tlb_entries_p0_d__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_31_addr = 5'h1a;
  assign tlb_entries_p0_d__T_31_data = tlb_entries_p0_d[tlb_entries_p0_d__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_32_addr = 5'h1b;
  assign tlb_entries_p0_d__T_32_data = tlb_entries_p0_d[tlb_entries_p0_d__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_33_addr = 5'h1c;
  assign tlb_entries_p0_d__T_33_data = tlb_entries_p0_d[tlb_entries_p0_d__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_34_addr = 5'h1d;
  assign tlb_entries_p0_d__T_34_data = tlb_entries_p0_d[tlb_entries_p0_d__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_35_addr = 5'h1e;
  assign tlb_entries_p0_d__T_35_data = tlb_entries_p0_d[tlb_entries_p0_d__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_36_addr = 5'h1f;
  assign tlb_entries_p0_d__T_36_data = tlb_entries_p0_d[tlb_entries_p0_d__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1546_addr = 5'h0;
  assign tlb_entries_p0_d__T_1546_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1547_addr = 5'h1;
  assign tlb_entries_p0_d__T_1547_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1548_addr = 5'h2;
  assign tlb_entries_p0_d__T_1548_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1549_addr = 5'h3;
  assign tlb_entries_p0_d__T_1549_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1550_addr = 5'h4;
  assign tlb_entries_p0_d__T_1550_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1551_addr = 5'h5;
  assign tlb_entries_p0_d__T_1551_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1552_addr = 5'h6;
  assign tlb_entries_p0_d__T_1552_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1553_addr = 5'h7;
  assign tlb_entries_p0_d__T_1553_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1554_addr = 5'h8;
  assign tlb_entries_p0_d__T_1554_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1555_addr = 5'h9;
  assign tlb_entries_p0_d__T_1555_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1556_addr = 5'ha;
  assign tlb_entries_p0_d__T_1556_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1557_addr = 5'hb;
  assign tlb_entries_p0_d__T_1557_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1558_addr = 5'hc;
  assign tlb_entries_p0_d__T_1558_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1559_addr = 5'hd;
  assign tlb_entries_p0_d__T_1559_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1560_addr = 5'he;
  assign tlb_entries_p0_d__T_1560_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1561_addr = 5'hf;
  assign tlb_entries_p0_d__T_1561_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1562_addr = 5'h10;
  assign tlb_entries_p0_d__T_1562_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1563_addr = 5'h11;
  assign tlb_entries_p0_d__T_1563_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1564_addr = 5'h12;
  assign tlb_entries_p0_d__T_1564_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1565_addr = 5'h13;
  assign tlb_entries_p0_d__T_1565_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1566_addr = 5'h14;
  assign tlb_entries_p0_d__T_1566_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1567_addr = 5'h15;
  assign tlb_entries_p0_d__T_1567_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1568_addr = 5'h16;
  assign tlb_entries_p0_d__T_1568_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1569_addr = 5'h17;
  assign tlb_entries_p0_d__T_1569_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1570_addr = 5'h18;
  assign tlb_entries_p0_d__T_1570_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1571_addr = 5'h19;
  assign tlb_entries_p0_d__T_1571_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1572_addr = 5'h1a;
  assign tlb_entries_p0_d__T_1572_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1573_addr = 5'h1b;
  assign tlb_entries_p0_d__T_1573_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1574_addr = 5'h1c;
  assign tlb_entries_p0_d__T_1574_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1575_addr = 5'h1d;
  assign tlb_entries_p0_d__T_1575_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1576_addr = 5'h1e;
  assign tlb_entries_p0_d__T_1576_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d__T_1577_addr = 5'h1f;
  assign tlb_entries_p0_d__T_1577_data = tlb_entries_p0_d[tlb_entries_p0_d__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p0_d_tlb_entry_ports_0_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p0_d_tlb_entry_ports_1_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p0_d_tlb_entry_ports_2_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p0_d_tlb_entry_ports_3_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p0_d_tlb_entry_ports_4_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p0_d_tlb_entry_ports_5_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p0_d_tlb_entry_ports_6_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p0_d_tlb_entry_ports_7_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p0_d_tlb_entry_ports_8_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p0_d_tlb_entry_ports_9_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p0_d_tlb_entry_ports_10_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p0_d_tlb_entry_ports_11_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p0_d_tlb_entry_ports_12_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p0_d_tlb_entry_ports_13_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p0_d_tlb_entry_ports_14_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p0_d_tlb_entry_ports_15_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p0_d_tlb_entry_ports_16_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p0_d_tlb_entry_ports_17_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p0_d_tlb_entry_ports_18_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p0_d_tlb_entry_ports_19_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p0_d_tlb_entry_ports_20_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p0_d_tlb_entry_ports_21_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p0_d_tlb_entry_ports_22_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p0_d_tlb_entry_ports_23_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p0_d_tlb_entry_ports_24_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p0_d_tlb_entry_ports_25_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p0_d_tlb_entry_ports_26_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p0_d_tlb_entry_ports_27_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p0_d_tlb_entry_ports_28_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p0_d_tlb_entry_ports_29_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p0_d_tlb_entry_ports_30_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p0_d_tlb_entry_ports_31_r_data = tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_d_tlb_entry_ports_0_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p0_d_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p0_d_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p0_d_tlb_entry_ports_1_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p0_d_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p0_d_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p0_d_tlb_entry_ports_2_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p0_d_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p0_d_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p0_d_tlb_entry_ports_3_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p0_d_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p0_d_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p0_d_tlb_entry_ports_4_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p0_d_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p0_d_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p0_d_tlb_entry_ports_5_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p0_d_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p0_d_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p0_d_tlb_entry_ports_6_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p0_d_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p0_d_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p0_d_tlb_entry_ports_7_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p0_d_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p0_d_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p0_d_tlb_entry_ports_8_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p0_d_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p0_d_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p0_d_tlb_entry_ports_9_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p0_d_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p0_d_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p0_d_tlb_entry_ports_10_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p0_d_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p0_d_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p0_d_tlb_entry_ports_11_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p0_d_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p0_d_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p0_d_tlb_entry_ports_12_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p0_d_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p0_d_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p0_d_tlb_entry_ports_13_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p0_d_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p0_d_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p0_d_tlb_entry_ports_14_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p0_d_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p0_d_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p0_d_tlb_entry_ports_15_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p0_d_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p0_d_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p0_d_tlb_entry_ports_16_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p0_d_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p0_d_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p0_d_tlb_entry_ports_17_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p0_d_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p0_d_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p0_d_tlb_entry_ports_18_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p0_d_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p0_d_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p0_d_tlb_entry_ports_19_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p0_d_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p0_d_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p0_d_tlb_entry_ports_20_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p0_d_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p0_d_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p0_d_tlb_entry_ports_21_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p0_d_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p0_d_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p0_d_tlb_entry_ports_22_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p0_d_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p0_d_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p0_d_tlb_entry_ports_23_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p0_d_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p0_d_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p0_d_tlb_entry_ports_24_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p0_d_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p0_d_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p0_d_tlb_entry_ports_25_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p0_d_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p0_d_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p0_d_tlb_entry_ports_26_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p0_d_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p0_d_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p0_d_tlb_entry_ports_27_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p0_d_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p0_d_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p0_d_tlb_entry_ports_28_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p0_d_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p0_d_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p0_d_tlb_entry_ports_29_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p0_d_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p0_d_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p0_d_tlb_entry_ports_30_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p0_d_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p0_d_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p0_d_tlb_entry_ports_31_w_data = io_wport_bits_entry_p0_d;
  assign tlb_entries_p0_d_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p0_d_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p0_d_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p0_v__T_5_addr = 5'h0;
  assign tlb_entries_p0_v__T_5_data = tlb_entries_p0_v[tlb_entries_p0_v__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_6_addr = 5'h1;
  assign tlb_entries_p0_v__T_6_data = tlb_entries_p0_v[tlb_entries_p0_v__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_7_addr = 5'h2;
  assign tlb_entries_p0_v__T_7_data = tlb_entries_p0_v[tlb_entries_p0_v__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_8_addr = 5'h3;
  assign tlb_entries_p0_v__T_8_data = tlb_entries_p0_v[tlb_entries_p0_v__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_9_addr = 5'h4;
  assign tlb_entries_p0_v__T_9_data = tlb_entries_p0_v[tlb_entries_p0_v__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_10_addr = 5'h5;
  assign tlb_entries_p0_v__T_10_data = tlb_entries_p0_v[tlb_entries_p0_v__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_11_addr = 5'h6;
  assign tlb_entries_p0_v__T_11_data = tlb_entries_p0_v[tlb_entries_p0_v__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_12_addr = 5'h7;
  assign tlb_entries_p0_v__T_12_data = tlb_entries_p0_v[tlb_entries_p0_v__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_13_addr = 5'h8;
  assign tlb_entries_p0_v__T_13_data = tlb_entries_p0_v[tlb_entries_p0_v__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_14_addr = 5'h9;
  assign tlb_entries_p0_v__T_14_data = tlb_entries_p0_v[tlb_entries_p0_v__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_15_addr = 5'ha;
  assign tlb_entries_p0_v__T_15_data = tlb_entries_p0_v[tlb_entries_p0_v__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_16_addr = 5'hb;
  assign tlb_entries_p0_v__T_16_data = tlb_entries_p0_v[tlb_entries_p0_v__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_17_addr = 5'hc;
  assign tlb_entries_p0_v__T_17_data = tlb_entries_p0_v[tlb_entries_p0_v__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_18_addr = 5'hd;
  assign tlb_entries_p0_v__T_18_data = tlb_entries_p0_v[tlb_entries_p0_v__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_19_addr = 5'he;
  assign tlb_entries_p0_v__T_19_data = tlb_entries_p0_v[tlb_entries_p0_v__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_20_addr = 5'hf;
  assign tlb_entries_p0_v__T_20_data = tlb_entries_p0_v[tlb_entries_p0_v__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_21_addr = 5'h10;
  assign tlb_entries_p0_v__T_21_data = tlb_entries_p0_v[tlb_entries_p0_v__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_22_addr = 5'h11;
  assign tlb_entries_p0_v__T_22_data = tlb_entries_p0_v[tlb_entries_p0_v__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_23_addr = 5'h12;
  assign tlb_entries_p0_v__T_23_data = tlb_entries_p0_v[tlb_entries_p0_v__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_24_addr = 5'h13;
  assign tlb_entries_p0_v__T_24_data = tlb_entries_p0_v[tlb_entries_p0_v__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_25_addr = 5'h14;
  assign tlb_entries_p0_v__T_25_data = tlb_entries_p0_v[tlb_entries_p0_v__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_26_addr = 5'h15;
  assign tlb_entries_p0_v__T_26_data = tlb_entries_p0_v[tlb_entries_p0_v__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_27_addr = 5'h16;
  assign tlb_entries_p0_v__T_27_data = tlb_entries_p0_v[tlb_entries_p0_v__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_28_addr = 5'h17;
  assign tlb_entries_p0_v__T_28_data = tlb_entries_p0_v[tlb_entries_p0_v__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_29_addr = 5'h18;
  assign tlb_entries_p0_v__T_29_data = tlb_entries_p0_v[tlb_entries_p0_v__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_30_addr = 5'h19;
  assign tlb_entries_p0_v__T_30_data = tlb_entries_p0_v[tlb_entries_p0_v__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_31_addr = 5'h1a;
  assign tlb_entries_p0_v__T_31_data = tlb_entries_p0_v[tlb_entries_p0_v__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_32_addr = 5'h1b;
  assign tlb_entries_p0_v__T_32_data = tlb_entries_p0_v[tlb_entries_p0_v__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_33_addr = 5'h1c;
  assign tlb_entries_p0_v__T_33_data = tlb_entries_p0_v[tlb_entries_p0_v__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_34_addr = 5'h1d;
  assign tlb_entries_p0_v__T_34_data = tlb_entries_p0_v[tlb_entries_p0_v__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_35_addr = 5'h1e;
  assign tlb_entries_p0_v__T_35_data = tlb_entries_p0_v[tlb_entries_p0_v__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_36_addr = 5'h1f;
  assign tlb_entries_p0_v__T_36_data = tlb_entries_p0_v[tlb_entries_p0_v__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1546_addr = 5'h0;
  assign tlb_entries_p0_v__T_1546_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1547_addr = 5'h1;
  assign tlb_entries_p0_v__T_1547_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1548_addr = 5'h2;
  assign tlb_entries_p0_v__T_1548_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1549_addr = 5'h3;
  assign tlb_entries_p0_v__T_1549_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1550_addr = 5'h4;
  assign tlb_entries_p0_v__T_1550_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1551_addr = 5'h5;
  assign tlb_entries_p0_v__T_1551_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1552_addr = 5'h6;
  assign tlb_entries_p0_v__T_1552_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1553_addr = 5'h7;
  assign tlb_entries_p0_v__T_1553_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1554_addr = 5'h8;
  assign tlb_entries_p0_v__T_1554_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1555_addr = 5'h9;
  assign tlb_entries_p0_v__T_1555_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1556_addr = 5'ha;
  assign tlb_entries_p0_v__T_1556_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1557_addr = 5'hb;
  assign tlb_entries_p0_v__T_1557_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1558_addr = 5'hc;
  assign tlb_entries_p0_v__T_1558_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1559_addr = 5'hd;
  assign tlb_entries_p0_v__T_1559_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1560_addr = 5'he;
  assign tlb_entries_p0_v__T_1560_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1561_addr = 5'hf;
  assign tlb_entries_p0_v__T_1561_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1562_addr = 5'h10;
  assign tlb_entries_p0_v__T_1562_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1563_addr = 5'h11;
  assign tlb_entries_p0_v__T_1563_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1564_addr = 5'h12;
  assign tlb_entries_p0_v__T_1564_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1565_addr = 5'h13;
  assign tlb_entries_p0_v__T_1565_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1566_addr = 5'h14;
  assign tlb_entries_p0_v__T_1566_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1567_addr = 5'h15;
  assign tlb_entries_p0_v__T_1567_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1568_addr = 5'h16;
  assign tlb_entries_p0_v__T_1568_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1569_addr = 5'h17;
  assign tlb_entries_p0_v__T_1569_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1570_addr = 5'h18;
  assign tlb_entries_p0_v__T_1570_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1571_addr = 5'h19;
  assign tlb_entries_p0_v__T_1571_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1572_addr = 5'h1a;
  assign tlb_entries_p0_v__T_1572_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1573_addr = 5'h1b;
  assign tlb_entries_p0_v__T_1573_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1574_addr = 5'h1c;
  assign tlb_entries_p0_v__T_1574_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1575_addr = 5'h1d;
  assign tlb_entries_p0_v__T_1575_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1576_addr = 5'h1e;
  assign tlb_entries_p0_v__T_1576_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v__T_1577_addr = 5'h1f;
  assign tlb_entries_p0_v__T_1577_data = tlb_entries_p0_v[tlb_entries_p0_v__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p0_v_tlb_entry_ports_0_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p0_v_tlb_entry_ports_1_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p0_v_tlb_entry_ports_2_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p0_v_tlb_entry_ports_3_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p0_v_tlb_entry_ports_4_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p0_v_tlb_entry_ports_5_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p0_v_tlb_entry_ports_6_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p0_v_tlb_entry_ports_7_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p0_v_tlb_entry_ports_8_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p0_v_tlb_entry_ports_9_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p0_v_tlb_entry_ports_10_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p0_v_tlb_entry_ports_11_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p0_v_tlb_entry_ports_12_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p0_v_tlb_entry_ports_13_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p0_v_tlb_entry_ports_14_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p0_v_tlb_entry_ports_15_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p0_v_tlb_entry_ports_16_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p0_v_tlb_entry_ports_17_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p0_v_tlb_entry_ports_18_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p0_v_tlb_entry_ports_19_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p0_v_tlb_entry_ports_20_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p0_v_tlb_entry_ports_21_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p0_v_tlb_entry_ports_22_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p0_v_tlb_entry_ports_23_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p0_v_tlb_entry_ports_24_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p0_v_tlb_entry_ports_25_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p0_v_tlb_entry_ports_26_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p0_v_tlb_entry_ports_27_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p0_v_tlb_entry_ports_28_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p0_v_tlb_entry_ports_29_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p0_v_tlb_entry_ports_30_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p0_v_tlb_entry_ports_31_r_data = tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p0_v_tlb_entry_ports_0_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p0_v_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p0_v_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p0_v_tlb_entry_ports_1_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p0_v_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p0_v_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p0_v_tlb_entry_ports_2_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p0_v_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p0_v_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p0_v_tlb_entry_ports_3_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p0_v_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p0_v_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p0_v_tlb_entry_ports_4_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p0_v_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p0_v_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p0_v_tlb_entry_ports_5_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p0_v_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p0_v_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p0_v_tlb_entry_ports_6_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p0_v_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p0_v_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p0_v_tlb_entry_ports_7_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p0_v_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p0_v_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p0_v_tlb_entry_ports_8_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p0_v_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p0_v_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p0_v_tlb_entry_ports_9_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p0_v_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p0_v_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p0_v_tlb_entry_ports_10_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p0_v_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p0_v_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p0_v_tlb_entry_ports_11_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p0_v_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p0_v_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p0_v_tlb_entry_ports_12_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p0_v_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p0_v_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p0_v_tlb_entry_ports_13_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p0_v_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p0_v_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p0_v_tlb_entry_ports_14_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p0_v_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p0_v_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p0_v_tlb_entry_ports_15_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p0_v_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p0_v_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p0_v_tlb_entry_ports_16_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p0_v_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p0_v_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p0_v_tlb_entry_ports_17_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p0_v_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p0_v_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p0_v_tlb_entry_ports_18_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p0_v_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p0_v_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p0_v_tlb_entry_ports_19_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p0_v_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p0_v_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p0_v_tlb_entry_ports_20_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p0_v_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p0_v_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p0_v_tlb_entry_ports_21_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p0_v_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p0_v_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p0_v_tlb_entry_ports_22_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p0_v_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p0_v_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p0_v_tlb_entry_ports_23_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p0_v_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p0_v_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p0_v_tlb_entry_ports_24_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p0_v_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p0_v_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p0_v_tlb_entry_ports_25_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p0_v_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p0_v_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p0_v_tlb_entry_ports_26_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p0_v_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p0_v_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p0_v_tlb_entry_ports_27_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p0_v_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p0_v_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p0_v_tlb_entry_ports_28_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p0_v_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p0_v_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p0_v_tlb_entry_ports_29_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p0_v_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p0_v_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p0_v_tlb_entry_ports_30_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p0_v_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p0_v_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p0_v_tlb_entry_ports_31_w_data = io_wport_bits_entry_p0_v;
  assign tlb_entries_p0_v_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p0_v_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p0_v_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p1_pfn__T_5_addr = 5'h0;
  assign tlb_entries_p1_pfn__T_5_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_6_addr = 5'h1;
  assign tlb_entries_p1_pfn__T_6_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_7_addr = 5'h2;
  assign tlb_entries_p1_pfn__T_7_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_8_addr = 5'h3;
  assign tlb_entries_p1_pfn__T_8_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_9_addr = 5'h4;
  assign tlb_entries_p1_pfn__T_9_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_10_addr = 5'h5;
  assign tlb_entries_p1_pfn__T_10_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_11_addr = 5'h6;
  assign tlb_entries_p1_pfn__T_11_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_12_addr = 5'h7;
  assign tlb_entries_p1_pfn__T_12_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_13_addr = 5'h8;
  assign tlb_entries_p1_pfn__T_13_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_14_addr = 5'h9;
  assign tlb_entries_p1_pfn__T_14_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_15_addr = 5'ha;
  assign tlb_entries_p1_pfn__T_15_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_16_addr = 5'hb;
  assign tlb_entries_p1_pfn__T_16_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_17_addr = 5'hc;
  assign tlb_entries_p1_pfn__T_17_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_18_addr = 5'hd;
  assign tlb_entries_p1_pfn__T_18_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_19_addr = 5'he;
  assign tlb_entries_p1_pfn__T_19_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_20_addr = 5'hf;
  assign tlb_entries_p1_pfn__T_20_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_21_addr = 5'h10;
  assign tlb_entries_p1_pfn__T_21_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_22_addr = 5'h11;
  assign tlb_entries_p1_pfn__T_22_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_23_addr = 5'h12;
  assign tlb_entries_p1_pfn__T_23_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_24_addr = 5'h13;
  assign tlb_entries_p1_pfn__T_24_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_25_addr = 5'h14;
  assign tlb_entries_p1_pfn__T_25_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_26_addr = 5'h15;
  assign tlb_entries_p1_pfn__T_26_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_27_addr = 5'h16;
  assign tlb_entries_p1_pfn__T_27_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_28_addr = 5'h17;
  assign tlb_entries_p1_pfn__T_28_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_29_addr = 5'h18;
  assign tlb_entries_p1_pfn__T_29_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_30_addr = 5'h19;
  assign tlb_entries_p1_pfn__T_30_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_31_addr = 5'h1a;
  assign tlb_entries_p1_pfn__T_31_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_32_addr = 5'h1b;
  assign tlb_entries_p1_pfn__T_32_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_33_addr = 5'h1c;
  assign tlb_entries_p1_pfn__T_33_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_34_addr = 5'h1d;
  assign tlb_entries_p1_pfn__T_34_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_35_addr = 5'h1e;
  assign tlb_entries_p1_pfn__T_35_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_36_addr = 5'h1f;
  assign tlb_entries_p1_pfn__T_36_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1546_addr = 5'h0;
  assign tlb_entries_p1_pfn__T_1546_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1547_addr = 5'h1;
  assign tlb_entries_p1_pfn__T_1547_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1548_addr = 5'h2;
  assign tlb_entries_p1_pfn__T_1548_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1549_addr = 5'h3;
  assign tlb_entries_p1_pfn__T_1549_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1550_addr = 5'h4;
  assign tlb_entries_p1_pfn__T_1550_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1551_addr = 5'h5;
  assign tlb_entries_p1_pfn__T_1551_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1552_addr = 5'h6;
  assign tlb_entries_p1_pfn__T_1552_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1553_addr = 5'h7;
  assign tlb_entries_p1_pfn__T_1553_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1554_addr = 5'h8;
  assign tlb_entries_p1_pfn__T_1554_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1555_addr = 5'h9;
  assign tlb_entries_p1_pfn__T_1555_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1556_addr = 5'ha;
  assign tlb_entries_p1_pfn__T_1556_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1557_addr = 5'hb;
  assign tlb_entries_p1_pfn__T_1557_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1558_addr = 5'hc;
  assign tlb_entries_p1_pfn__T_1558_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1559_addr = 5'hd;
  assign tlb_entries_p1_pfn__T_1559_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1560_addr = 5'he;
  assign tlb_entries_p1_pfn__T_1560_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1561_addr = 5'hf;
  assign tlb_entries_p1_pfn__T_1561_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1562_addr = 5'h10;
  assign tlb_entries_p1_pfn__T_1562_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1563_addr = 5'h11;
  assign tlb_entries_p1_pfn__T_1563_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1564_addr = 5'h12;
  assign tlb_entries_p1_pfn__T_1564_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1565_addr = 5'h13;
  assign tlb_entries_p1_pfn__T_1565_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1566_addr = 5'h14;
  assign tlb_entries_p1_pfn__T_1566_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1567_addr = 5'h15;
  assign tlb_entries_p1_pfn__T_1567_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1568_addr = 5'h16;
  assign tlb_entries_p1_pfn__T_1568_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1569_addr = 5'h17;
  assign tlb_entries_p1_pfn__T_1569_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1570_addr = 5'h18;
  assign tlb_entries_p1_pfn__T_1570_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1571_addr = 5'h19;
  assign tlb_entries_p1_pfn__T_1571_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1572_addr = 5'h1a;
  assign tlb_entries_p1_pfn__T_1572_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1573_addr = 5'h1b;
  assign tlb_entries_p1_pfn__T_1573_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1574_addr = 5'h1c;
  assign tlb_entries_p1_pfn__T_1574_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1575_addr = 5'h1d;
  assign tlb_entries_p1_pfn__T_1575_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1576_addr = 5'h1e;
  assign tlb_entries_p1_pfn__T_1576_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn__T_1577_addr = 5'h1f;
  assign tlb_entries_p1_pfn__T_1577_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p1_pfn_tlb_entry_ports_0_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p1_pfn_tlb_entry_ports_1_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p1_pfn_tlb_entry_ports_2_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p1_pfn_tlb_entry_ports_3_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p1_pfn_tlb_entry_ports_4_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p1_pfn_tlb_entry_ports_5_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p1_pfn_tlb_entry_ports_6_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p1_pfn_tlb_entry_ports_7_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p1_pfn_tlb_entry_ports_8_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p1_pfn_tlb_entry_ports_9_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p1_pfn_tlb_entry_ports_10_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p1_pfn_tlb_entry_ports_11_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p1_pfn_tlb_entry_ports_12_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p1_pfn_tlb_entry_ports_13_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p1_pfn_tlb_entry_ports_14_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p1_pfn_tlb_entry_ports_15_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p1_pfn_tlb_entry_ports_16_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p1_pfn_tlb_entry_ports_17_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p1_pfn_tlb_entry_ports_18_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p1_pfn_tlb_entry_ports_19_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p1_pfn_tlb_entry_ports_20_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p1_pfn_tlb_entry_ports_21_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p1_pfn_tlb_entry_ports_22_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p1_pfn_tlb_entry_ports_23_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p1_pfn_tlb_entry_ports_24_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p1_pfn_tlb_entry_ports_25_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p1_pfn_tlb_entry_ports_26_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p1_pfn_tlb_entry_ports_27_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p1_pfn_tlb_entry_ports_28_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p1_pfn_tlb_entry_ports_29_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p1_pfn_tlb_entry_ports_30_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p1_pfn_tlb_entry_ports_31_r_data = tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_pfn_tlb_entry_ports_0_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p1_pfn_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p1_pfn_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p1_pfn_tlb_entry_ports_1_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p1_pfn_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p1_pfn_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p1_pfn_tlb_entry_ports_2_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p1_pfn_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p1_pfn_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p1_pfn_tlb_entry_ports_3_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p1_pfn_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p1_pfn_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p1_pfn_tlb_entry_ports_4_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p1_pfn_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p1_pfn_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p1_pfn_tlb_entry_ports_5_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p1_pfn_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p1_pfn_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p1_pfn_tlb_entry_ports_6_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p1_pfn_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p1_pfn_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p1_pfn_tlb_entry_ports_7_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p1_pfn_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p1_pfn_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p1_pfn_tlb_entry_ports_8_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p1_pfn_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p1_pfn_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p1_pfn_tlb_entry_ports_9_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p1_pfn_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p1_pfn_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p1_pfn_tlb_entry_ports_10_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p1_pfn_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p1_pfn_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p1_pfn_tlb_entry_ports_11_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p1_pfn_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p1_pfn_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p1_pfn_tlb_entry_ports_12_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p1_pfn_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p1_pfn_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p1_pfn_tlb_entry_ports_13_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p1_pfn_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p1_pfn_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p1_pfn_tlb_entry_ports_14_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p1_pfn_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p1_pfn_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p1_pfn_tlb_entry_ports_15_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p1_pfn_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p1_pfn_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p1_pfn_tlb_entry_ports_16_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p1_pfn_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p1_pfn_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p1_pfn_tlb_entry_ports_17_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p1_pfn_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p1_pfn_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p1_pfn_tlb_entry_ports_18_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p1_pfn_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p1_pfn_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p1_pfn_tlb_entry_ports_19_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p1_pfn_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p1_pfn_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p1_pfn_tlb_entry_ports_20_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p1_pfn_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p1_pfn_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p1_pfn_tlb_entry_ports_21_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p1_pfn_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p1_pfn_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p1_pfn_tlb_entry_ports_22_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p1_pfn_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p1_pfn_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p1_pfn_tlb_entry_ports_23_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p1_pfn_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p1_pfn_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p1_pfn_tlb_entry_ports_24_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p1_pfn_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p1_pfn_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p1_pfn_tlb_entry_ports_25_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p1_pfn_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p1_pfn_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p1_pfn_tlb_entry_ports_26_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p1_pfn_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p1_pfn_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p1_pfn_tlb_entry_ports_27_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p1_pfn_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p1_pfn_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p1_pfn_tlb_entry_ports_28_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p1_pfn_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p1_pfn_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p1_pfn_tlb_entry_ports_29_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p1_pfn_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p1_pfn_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p1_pfn_tlb_entry_ports_30_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p1_pfn_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p1_pfn_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p1_pfn_tlb_entry_ports_31_w_data = io_wport_bits_entry_p1_pfn;
  assign tlb_entries_p1_pfn_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p1_pfn_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p1_pfn_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p1_c__T_5_addr = 5'h0;
  assign tlb_entries_p1_c__T_5_data = tlb_entries_p1_c[tlb_entries_p1_c__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_6_addr = 5'h1;
  assign tlb_entries_p1_c__T_6_data = tlb_entries_p1_c[tlb_entries_p1_c__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_7_addr = 5'h2;
  assign tlb_entries_p1_c__T_7_data = tlb_entries_p1_c[tlb_entries_p1_c__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_8_addr = 5'h3;
  assign tlb_entries_p1_c__T_8_data = tlb_entries_p1_c[tlb_entries_p1_c__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_9_addr = 5'h4;
  assign tlb_entries_p1_c__T_9_data = tlb_entries_p1_c[tlb_entries_p1_c__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_10_addr = 5'h5;
  assign tlb_entries_p1_c__T_10_data = tlb_entries_p1_c[tlb_entries_p1_c__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_11_addr = 5'h6;
  assign tlb_entries_p1_c__T_11_data = tlb_entries_p1_c[tlb_entries_p1_c__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_12_addr = 5'h7;
  assign tlb_entries_p1_c__T_12_data = tlb_entries_p1_c[tlb_entries_p1_c__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_13_addr = 5'h8;
  assign tlb_entries_p1_c__T_13_data = tlb_entries_p1_c[tlb_entries_p1_c__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_14_addr = 5'h9;
  assign tlb_entries_p1_c__T_14_data = tlb_entries_p1_c[tlb_entries_p1_c__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_15_addr = 5'ha;
  assign tlb_entries_p1_c__T_15_data = tlb_entries_p1_c[tlb_entries_p1_c__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_16_addr = 5'hb;
  assign tlb_entries_p1_c__T_16_data = tlb_entries_p1_c[tlb_entries_p1_c__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_17_addr = 5'hc;
  assign tlb_entries_p1_c__T_17_data = tlb_entries_p1_c[tlb_entries_p1_c__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_18_addr = 5'hd;
  assign tlb_entries_p1_c__T_18_data = tlb_entries_p1_c[tlb_entries_p1_c__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_19_addr = 5'he;
  assign tlb_entries_p1_c__T_19_data = tlb_entries_p1_c[tlb_entries_p1_c__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_20_addr = 5'hf;
  assign tlb_entries_p1_c__T_20_data = tlb_entries_p1_c[tlb_entries_p1_c__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_21_addr = 5'h10;
  assign tlb_entries_p1_c__T_21_data = tlb_entries_p1_c[tlb_entries_p1_c__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_22_addr = 5'h11;
  assign tlb_entries_p1_c__T_22_data = tlb_entries_p1_c[tlb_entries_p1_c__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_23_addr = 5'h12;
  assign tlb_entries_p1_c__T_23_data = tlb_entries_p1_c[tlb_entries_p1_c__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_24_addr = 5'h13;
  assign tlb_entries_p1_c__T_24_data = tlb_entries_p1_c[tlb_entries_p1_c__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_25_addr = 5'h14;
  assign tlb_entries_p1_c__T_25_data = tlb_entries_p1_c[tlb_entries_p1_c__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_26_addr = 5'h15;
  assign tlb_entries_p1_c__T_26_data = tlb_entries_p1_c[tlb_entries_p1_c__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_27_addr = 5'h16;
  assign tlb_entries_p1_c__T_27_data = tlb_entries_p1_c[tlb_entries_p1_c__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_28_addr = 5'h17;
  assign tlb_entries_p1_c__T_28_data = tlb_entries_p1_c[tlb_entries_p1_c__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_29_addr = 5'h18;
  assign tlb_entries_p1_c__T_29_data = tlb_entries_p1_c[tlb_entries_p1_c__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_30_addr = 5'h19;
  assign tlb_entries_p1_c__T_30_data = tlb_entries_p1_c[tlb_entries_p1_c__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_31_addr = 5'h1a;
  assign tlb_entries_p1_c__T_31_data = tlb_entries_p1_c[tlb_entries_p1_c__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_32_addr = 5'h1b;
  assign tlb_entries_p1_c__T_32_data = tlb_entries_p1_c[tlb_entries_p1_c__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_33_addr = 5'h1c;
  assign tlb_entries_p1_c__T_33_data = tlb_entries_p1_c[tlb_entries_p1_c__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_34_addr = 5'h1d;
  assign tlb_entries_p1_c__T_34_data = tlb_entries_p1_c[tlb_entries_p1_c__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_35_addr = 5'h1e;
  assign tlb_entries_p1_c__T_35_data = tlb_entries_p1_c[tlb_entries_p1_c__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_36_addr = 5'h1f;
  assign tlb_entries_p1_c__T_36_data = tlb_entries_p1_c[tlb_entries_p1_c__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1546_addr = 5'h0;
  assign tlb_entries_p1_c__T_1546_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1547_addr = 5'h1;
  assign tlb_entries_p1_c__T_1547_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1548_addr = 5'h2;
  assign tlb_entries_p1_c__T_1548_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1549_addr = 5'h3;
  assign tlb_entries_p1_c__T_1549_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1550_addr = 5'h4;
  assign tlb_entries_p1_c__T_1550_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1551_addr = 5'h5;
  assign tlb_entries_p1_c__T_1551_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1552_addr = 5'h6;
  assign tlb_entries_p1_c__T_1552_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1553_addr = 5'h7;
  assign tlb_entries_p1_c__T_1553_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1554_addr = 5'h8;
  assign tlb_entries_p1_c__T_1554_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1555_addr = 5'h9;
  assign tlb_entries_p1_c__T_1555_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1556_addr = 5'ha;
  assign tlb_entries_p1_c__T_1556_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1557_addr = 5'hb;
  assign tlb_entries_p1_c__T_1557_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1558_addr = 5'hc;
  assign tlb_entries_p1_c__T_1558_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1559_addr = 5'hd;
  assign tlb_entries_p1_c__T_1559_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1560_addr = 5'he;
  assign tlb_entries_p1_c__T_1560_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1561_addr = 5'hf;
  assign tlb_entries_p1_c__T_1561_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1562_addr = 5'h10;
  assign tlb_entries_p1_c__T_1562_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1563_addr = 5'h11;
  assign tlb_entries_p1_c__T_1563_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1564_addr = 5'h12;
  assign tlb_entries_p1_c__T_1564_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1565_addr = 5'h13;
  assign tlb_entries_p1_c__T_1565_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1566_addr = 5'h14;
  assign tlb_entries_p1_c__T_1566_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1567_addr = 5'h15;
  assign tlb_entries_p1_c__T_1567_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1568_addr = 5'h16;
  assign tlb_entries_p1_c__T_1568_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1569_addr = 5'h17;
  assign tlb_entries_p1_c__T_1569_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1570_addr = 5'h18;
  assign tlb_entries_p1_c__T_1570_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1571_addr = 5'h19;
  assign tlb_entries_p1_c__T_1571_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1572_addr = 5'h1a;
  assign tlb_entries_p1_c__T_1572_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1573_addr = 5'h1b;
  assign tlb_entries_p1_c__T_1573_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1574_addr = 5'h1c;
  assign tlb_entries_p1_c__T_1574_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1575_addr = 5'h1d;
  assign tlb_entries_p1_c__T_1575_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1576_addr = 5'h1e;
  assign tlb_entries_p1_c__T_1576_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c__T_1577_addr = 5'h1f;
  assign tlb_entries_p1_c__T_1577_data = tlb_entries_p1_c[tlb_entries_p1_c__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p1_c_tlb_entry_ports_0_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p1_c_tlb_entry_ports_1_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p1_c_tlb_entry_ports_2_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p1_c_tlb_entry_ports_3_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p1_c_tlb_entry_ports_4_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p1_c_tlb_entry_ports_5_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p1_c_tlb_entry_ports_6_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p1_c_tlb_entry_ports_7_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p1_c_tlb_entry_ports_8_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p1_c_tlb_entry_ports_9_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p1_c_tlb_entry_ports_10_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p1_c_tlb_entry_ports_11_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p1_c_tlb_entry_ports_12_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p1_c_tlb_entry_ports_13_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p1_c_tlb_entry_ports_14_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p1_c_tlb_entry_ports_15_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p1_c_tlb_entry_ports_16_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p1_c_tlb_entry_ports_17_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p1_c_tlb_entry_ports_18_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p1_c_tlb_entry_ports_19_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p1_c_tlb_entry_ports_20_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p1_c_tlb_entry_ports_21_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p1_c_tlb_entry_ports_22_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p1_c_tlb_entry_ports_23_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p1_c_tlb_entry_ports_24_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p1_c_tlb_entry_ports_25_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p1_c_tlb_entry_ports_26_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p1_c_tlb_entry_ports_27_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p1_c_tlb_entry_ports_28_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p1_c_tlb_entry_ports_29_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p1_c_tlb_entry_ports_30_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p1_c_tlb_entry_ports_31_r_data = tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_c_tlb_entry_ports_0_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p1_c_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p1_c_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p1_c_tlb_entry_ports_1_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p1_c_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p1_c_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p1_c_tlb_entry_ports_2_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p1_c_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p1_c_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p1_c_tlb_entry_ports_3_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p1_c_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p1_c_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p1_c_tlb_entry_ports_4_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p1_c_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p1_c_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p1_c_tlb_entry_ports_5_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p1_c_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p1_c_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p1_c_tlb_entry_ports_6_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p1_c_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p1_c_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p1_c_tlb_entry_ports_7_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p1_c_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p1_c_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p1_c_tlb_entry_ports_8_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p1_c_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p1_c_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p1_c_tlb_entry_ports_9_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p1_c_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p1_c_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p1_c_tlb_entry_ports_10_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p1_c_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p1_c_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p1_c_tlb_entry_ports_11_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p1_c_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p1_c_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p1_c_tlb_entry_ports_12_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p1_c_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p1_c_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p1_c_tlb_entry_ports_13_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p1_c_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p1_c_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p1_c_tlb_entry_ports_14_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p1_c_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p1_c_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p1_c_tlb_entry_ports_15_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p1_c_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p1_c_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p1_c_tlb_entry_ports_16_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p1_c_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p1_c_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p1_c_tlb_entry_ports_17_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p1_c_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p1_c_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p1_c_tlb_entry_ports_18_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p1_c_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p1_c_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p1_c_tlb_entry_ports_19_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p1_c_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p1_c_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p1_c_tlb_entry_ports_20_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p1_c_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p1_c_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p1_c_tlb_entry_ports_21_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p1_c_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p1_c_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p1_c_tlb_entry_ports_22_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p1_c_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p1_c_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p1_c_tlb_entry_ports_23_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p1_c_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p1_c_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p1_c_tlb_entry_ports_24_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p1_c_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p1_c_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p1_c_tlb_entry_ports_25_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p1_c_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p1_c_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p1_c_tlb_entry_ports_26_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p1_c_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p1_c_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p1_c_tlb_entry_ports_27_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p1_c_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p1_c_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p1_c_tlb_entry_ports_28_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p1_c_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p1_c_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p1_c_tlb_entry_ports_29_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p1_c_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p1_c_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p1_c_tlb_entry_ports_30_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p1_c_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p1_c_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p1_c_tlb_entry_ports_31_w_data = io_wport_bits_entry_p1_c;
  assign tlb_entries_p1_c_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p1_c_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p1_c_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p1_d__T_5_addr = 5'h0;
  assign tlb_entries_p1_d__T_5_data = tlb_entries_p1_d[tlb_entries_p1_d__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_6_addr = 5'h1;
  assign tlb_entries_p1_d__T_6_data = tlb_entries_p1_d[tlb_entries_p1_d__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_7_addr = 5'h2;
  assign tlb_entries_p1_d__T_7_data = tlb_entries_p1_d[tlb_entries_p1_d__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_8_addr = 5'h3;
  assign tlb_entries_p1_d__T_8_data = tlb_entries_p1_d[tlb_entries_p1_d__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_9_addr = 5'h4;
  assign tlb_entries_p1_d__T_9_data = tlb_entries_p1_d[tlb_entries_p1_d__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_10_addr = 5'h5;
  assign tlb_entries_p1_d__T_10_data = tlb_entries_p1_d[tlb_entries_p1_d__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_11_addr = 5'h6;
  assign tlb_entries_p1_d__T_11_data = tlb_entries_p1_d[tlb_entries_p1_d__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_12_addr = 5'h7;
  assign tlb_entries_p1_d__T_12_data = tlb_entries_p1_d[tlb_entries_p1_d__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_13_addr = 5'h8;
  assign tlb_entries_p1_d__T_13_data = tlb_entries_p1_d[tlb_entries_p1_d__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_14_addr = 5'h9;
  assign tlb_entries_p1_d__T_14_data = tlb_entries_p1_d[tlb_entries_p1_d__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_15_addr = 5'ha;
  assign tlb_entries_p1_d__T_15_data = tlb_entries_p1_d[tlb_entries_p1_d__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_16_addr = 5'hb;
  assign tlb_entries_p1_d__T_16_data = tlb_entries_p1_d[tlb_entries_p1_d__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_17_addr = 5'hc;
  assign tlb_entries_p1_d__T_17_data = tlb_entries_p1_d[tlb_entries_p1_d__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_18_addr = 5'hd;
  assign tlb_entries_p1_d__T_18_data = tlb_entries_p1_d[tlb_entries_p1_d__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_19_addr = 5'he;
  assign tlb_entries_p1_d__T_19_data = tlb_entries_p1_d[tlb_entries_p1_d__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_20_addr = 5'hf;
  assign tlb_entries_p1_d__T_20_data = tlb_entries_p1_d[tlb_entries_p1_d__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_21_addr = 5'h10;
  assign tlb_entries_p1_d__T_21_data = tlb_entries_p1_d[tlb_entries_p1_d__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_22_addr = 5'h11;
  assign tlb_entries_p1_d__T_22_data = tlb_entries_p1_d[tlb_entries_p1_d__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_23_addr = 5'h12;
  assign tlb_entries_p1_d__T_23_data = tlb_entries_p1_d[tlb_entries_p1_d__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_24_addr = 5'h13;
  assign tlb_entries_p1_d__T_24_data = tlb_entries_p1_d[tlb_entries_p1_d__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_25_addr = 5'h14;
  assign tlb_entries_p1_d__T_25_data = tlb_entries_p1_d[tlb_entries_p1_d__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_26_addr = 5'h15;
  assign tlb_entries_p1_d__T_26_data = tlb_entries_p1_d[tlb_entries_p1_d__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_27_addr = 5'h16;
  assign tlb_entries_p1_d__T_27_data = tlb_entries_p1_d[tlb_entries_p1_d__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_28_addr = 5'h17;
  assign tlb_entries_p1_d__T_28_data = tlb_entries_p1_d[tlb_entries_p1_d__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_29_addr = 5'h18;
  assign tlb_entries_p1_d__T_29_data = tlb_entries_p1_d[tlb_entries_p1_d__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_30_addr = 5'h19;
  assign tlb_entries_p1_d__T_30_data = tlb_entries_p1_d[tlb_entries_p1_d__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_31_addr = 5'h1a;
  assign tlb_entries_p1_d__T_31_data = tlb_entries_p1_d[tlb_entries_p1_d__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_32_addr = 5'h1b;
  assign tlb_entries_p1_d__T_32_data = tlb_entries_p1_d[tlb_entries_p1_d__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_33_addr = 5'h1c;
  assign tlb_entries_p1_d__T_33_data = tlb_entries_p1_d[tlb_entries_p1_d__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_34_addr = 5'h1d;
  assign tlb_entries_p1_d__T_34_data = tlb_entries_p1_d[tlb_entries_p1_d__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_35_addr = 5'h1e;
  assign tlb_entries_p1_d__T_35_data = tlb_entries_p1_d[tlb_entries_p1_d__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_36_addr = 5'h1f;
  assign tlb_entries_p1_d__T_36_data = tlb_entries_p1_d[tlb_entries_p1_d__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1546_addr = 5'h0;
  assign tlb_entries_p1_d__T_1546_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1547_addr = 5'h1;
  assign tlb_entries_p1_d__T_1547_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1548_addr = 5'h2;
  assign tlb_entries_p1_d__T_1548_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1549_addr = 5'h3;
  assign tlb_entries_p1_d__T_1549_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1550_addr = 5'h4;
  assign tlb_entries_p1_d__T_1550_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1551_addr = 5'h5;
  assign tlb_entries_p1_d__T_1551_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1552_addr = 5'h6;
  assign tlb_entries_p1_d__T_1552_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1553_addr = 5'h7;
  assign tlb_entries_p1_d__T_1553_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1554_addr = 5'h8;
  assign tlb_entries_p1_d__T_1554_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1555_addr = 5'h9;
  assign tlb_entries_p1_d__T_1555_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1556_addr = 5'ha;
  assign tlb_entries_p1_d__T_1556_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1557_addr = 5'hb;
  assign tlb_entries_p1_d__T_1557_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1558_addr = 5'hc;
  assign tlb_entries_p1_d__T_1558_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1559_addr = 5'hd;
  assign tlb_entries_p1_d__T_1559_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1560_addr = 5'he;
  assign tlb_entries_p1_d__T_1560_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1561_addr = 5'hf;
  assign tlb_entries_p1_d__T_1561_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1562_addr = 5'h10;
  assign tlb_entries_p1_d__T_1562_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1563_addr = 5'h11;
  assign tlb_entries_p1_d__T_1563_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1564_addr = 5'h12;
  assign tlb_entries_p1_d__T_1564_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1565_addr = 5'h13;
  assign tlb_entries_p1_d__T_1565_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1566_addr = 5'h14;
  assign tlb_entries_p1_d__T_1566_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1567_addr = 5'h15;
  assign tlb_entries_p1_d__T_1567_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1568_addr = 5'h16;
  assign tlb_entries_p1_d__T_1568_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1569_addr = 5'h17;
  assign tlb_entries_p1_d__T_1569_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1570_addr = 5'h18;
  assign tlb_entries_p1_d__T_1570_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1571_addr = 5'h19;
  assign tlb_entries_p1_d__T_1571_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1572_addr = 5'h1a;
  assign tlb_entries_p1_d__T_1572_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1573_addr = 5'h1b;
  assign tlb_entries_p1_d__T_1573_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1574_addr = 5'h1c;
  assign tlb_entries_p1_d__T_1574_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1575_addr = 5'h1d;
  assign tlb_entries_p1_d__T_1575_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1576_addr = 5'h1e;
  assign tlb_entries_p1_d__T_1576_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d__T_1577_addr = 5'h1f;
  assign tlb_entries_p1_d__T_1577_data = tlb_entries_p1_d[tlb_entries_p1_d__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p1_d_tlb_entry_ports_0_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p1_d_tlb_entry_ports_1_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p1_d_tlb_entry_ports_2_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p1_d_tlb_entry_ports_3_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p1_d_tlb_entry_ports_4_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p1_d_tlb_entry_ports_5_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p1_d_tlb_entry_ports_6_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p1_d_tlb_entry_ports_7_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p1_d_tlb_entry_ports_8_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p1_d_tlb_entry_ports_9_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p1_d_tlb_entry_ports_10_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p1_d_tlb_entry_ports_11_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p1_d_tlb_entry_ports_12_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p1_d_tlb_entry_ports_13_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p1_d_tlb_entry_ports_14_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p1_d_tlb_entry_ports_15_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p1_d_tlb_entry_ports_16_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p1_d_tlb_entry_ports_17_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p1_d_tlb_entry_ports_18_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p1_d_tlb_entry_ports_19_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p1_d_tlb_entry_ports_20_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p1_d_tlb_entry_ports_21_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p1_d_tlb_entry_ports_22_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p1_d_tlb_entry_ports_23_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p1_d_tlb_entry_ports_24_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p1_d_tlb_entry_ports_25_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p1_d_tlb_entry_ports_26_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p1_d_tlb_entry_ports_27_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p1_d_tlb_entry_ports_28_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p1_d_tlb_entry_ports_29_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p1_d_tlb_entry_ports_30_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p1_d_tlb_entry_ports_31_r_data = tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_d_tlb_entry_ports_0_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p1_d_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p1_d_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p1_d_tlb_entry_ports_1_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p1_d_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p1_d_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p1_d_tlb_entry_ports_2_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p1_d_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p1_d_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p1_d_tlb_entry_ports_3_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p1_d_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p1_d_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p1_d_tlb_entry_ports_4_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p1_d_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p1_d_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p1_d_tlb_entry_ports_5_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p1_d_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p1_d_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p1_d_tlb_entry_ports_6_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p1_d_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p1_d_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p1_d_tlb_entry_ports_7_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p1_d_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p1_d_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p1_d_tlb_entry_ports_8_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p1_d_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p1_d_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p1_d_tlb_entry_ports_9_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p1_d_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p1_d_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p1_d_tlb_entry_ports_10_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p1_d_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p1_d_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p1_d_tlb_entry_ports_11_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p1_d_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p1_d_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p1_d_tlb_entry_ports_12_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p1_d_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p1_d_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p1_d_tlb_entry_ports_13_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p1_d_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p1_d_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p1_d_tlb_entry_ports_14_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p1_d_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p1_d_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p1_d_tlb_entry_ports_15_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p1_d_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p1_d_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p1_d_tlb_entry_ports_16_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p1_d_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p1_d_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p1_d_tlb_entry_ports_17_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p1_d_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p1_d_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p1_d_tlb_entry_ports_18_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p1_d_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p1_d_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p1_d_tlb_entry_ports_19_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p1_d_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p1_d_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p1_d_tlb_entry_ports_20_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p1_d_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p1_d_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p1_d_tlb_entry_ports_21_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p1_d_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p1_d_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p1_d_tlb_entry_ports_22_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p1_d_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p1_d_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p1_d_tlb_entry_ports_23_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p1_d_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p1_d_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p1_d_tlb_entry_ports_24_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p1_d_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p1_d_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p1_d_tlb_entry_ports_25_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p1_d_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p1_d_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p1_d_tlb_entry_ports_26_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p1_d_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p1_d_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p1_d_tlb_entry_ports_27_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p1_d_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p1_d_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p1_d_tlb_entry_ports_28_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p1_d_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p1_d_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p1_d_tlb_entry_ports_29_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p1_d_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p1_d_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p1_d_tlb_entry_ports_30_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p1_d_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p1_d_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p1_d_tlb_entry_ports_31_w_data = io_wport_bits_entry_p1_d;
  assign tlb_entries_p1_d_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p1_d_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p1_d_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign tlb_entries_p1_v__T_5_addr = 5'h0;
  assign tlb_entries_p1_v__T_5_data = tlb_entries_p1_v[tlb_entries_p1_v__T_5_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_6_addr = 5'h1;
  assign tlb_entries_p1_v__T_6_data = tlb_entries_p1_v[tlb_entries_p1_v__T_6_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_7_addr = 5'h2;
  assign tlb_entries_p1_v__T_7_data = tlb_entries_p1_v[tlb_entries_p1_v__T_7_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_8_addr = 5'h3;
  assign tlb_entries_p1_v__T_8_data = tlb_entries_p1_v[tlb_entries_p1_v__T_8_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_9_addr = 5'h4;
  assign tlb_entries_p1_v__T_9_data = tlb_entries_p1_v[tlb_entries_p1_v__T_9_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_10_addr = 5'h5;
  assign tlb_entries_p1_v__T_10_data = tlb_entries_p1_v[tlb_entries_p1_v__T_10_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_11_addr = 5'h6;
  assign tlb_entries_p1_v__T_11_data = tlb_entries_p1_v[tlb_entries_p1_v__T_11_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_12_addr = 5'h7;
  assign tlb_entries_p1_v__T_12_data = tlb_entries_p1_v[tlb_entries_p1_v__T_12_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_13_addr = 5'h8;
  assign tlb_entries_p1_v__T_13_data = tlb_entries_p1_v[tlb_entries_p1_v__T_13_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_14_addr = 5'h9;
  assign tlb_entries_p1_v__T_14_data = tlb_entries_p1_v[tlb_entries_p1_v__T_14_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_15_addr = 5'ha;
  assign tlb_entries_p1_v__T_15_data = tlb_entries_p1_v[tlb_entries_p1_v__T_15_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_16_addr = 5'hb;
  assign tlb_entries_p1_v__T_16_data = tlb_entries_p1_v[tlb_entries_p1_v__T_16_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_17_addr = 5'hc;
  assign tlb_entries_p1_v__T_17_data = tlb_entries_p1_v[tlb_entries_p1_v__T_17_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_18_addr = 5'hd;
  assign tlb_entries_p1_v__T_18_data = tlb_entries_p1_v[tlb_entries_p1_v__T_18_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_19_addr = 5'he;
  assign tlb_entries_p1_v__T_19_data = tlb_entries_p1_v[tlb_entries_p1_v__T_19_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_20_addr = 5'hf;
  assign tlb_entries_p1_v__T_20_data = tlb_entries_p1_v[tlb_entries_p1_v__T_20_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_21_addr = 5'h10;
  assign tlb_entries_p1_v__T_21_data = tlb_entries_p1_v[tlb_entries_p1_v__T_21_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_22_addr = 5'h11;
  assign tlb_entries_p1_v__T_22_data = tlb_entries_p1_v[tlb_entries_p1_v__T_22_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_23_addr = 5'h12;
  assign tlb_entries_p1_v__T_23_data = tlb_entries_p1_v[tlb_entries_p1_v__T_23_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_24_addr = 5'h13;
  assign tlb_entries_p1_v__T_24_data = tlb_entries_p1_v[tlb_entries_p1_v__T_24_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_25_addr = 5'h14;
  assign tlb_entries_p1_v__T_25_data = tlb_entries_p1_v[tlb_entries_p1_v__T_25_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_26_addr = 5'h15;
  assign tlb_entries_p1_v__T_26_data = tlb_entries_p1_v[tlb_entries_p1_v__T_26_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_27_addr = 5'h16;
  assign tlb_entries_p1_v__T_27_data = tlb_entries_p1_v[tlb_entries_p1_v__T_27_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_28_addr = 5'h17;
  assign tlb_entries_p1_v__T_28_data = tlb_entries_p1_v[tlb_entries_p1_v__T_28_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_29_addr = 5'h18;
  assign tlb_entries_p1_v__T_29_data = tlb_entries_p1_v[tlb_entries_p1_v__T_29_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_30_addr = 5'h19;
  assign tlb_entries_p1_v__T_30_data = tlb_entries_p1_v[tlb_entries_p1_v__T_30_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_31_addr = 5'h1a;
  assign tlb_entries_p1_v__T_31_data = tlb_entries_p1_v[tlb_entries_p1_v__T_31_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_32_addr = 5'h1b;
  assign tlb_entries_p1_v__T_32_data = tlb_entries_p1_v[tlb_entries_p1_v__T_32_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_33_addr = 5'h1c;
  assign tlb_entries_p1_v__T_33_data = tlb_entries_p1_v[tlb_entries_p1_v__T_33_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_34_addr = 5'h1d;
  assign tlb_entries_p1_v__T_34_data = tlb_entries_p1_v[tlb_entries_p1_v__T_34_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_35_addr = 5'h1e;
  assign tlb_entries_p1_v__T_35_data = tlb_entries_p1_v[tlb_entries_p1_v__T_35_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_36_addr = 5'h1f;
  assign tlb_entries_p1_v__T_36_data = tlb_entries_p1_v[tlb_entries_p1_v__T_36_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1546_addr = 5'h0;
  assign tlb_entries_p1_v__T_1546_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1546_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1547_addr = 5'h1;
  assign tlb_entries_p1_v__T_1547_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1547_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1548_addr = 5'h2;
  assign tlb_entries_p1_v__T_1548_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1548_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1549_addr = 5'h3;
  assign tlb_entries_p1_v__T_1549_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1549_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1550_addr = 5'h4;
  assign tlb_entries_p1_v__T_1550_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1550_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1551_addr = 5'h5;
  assign tlb_entries_p1_v__T_1551_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1551_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1552_addr = 5'h6;
  assign tlb_entries_p1_v__T_1552_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1552_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1553_addr = 5'h7;
  assign tlb_entries_p1_v__T_1553_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1553_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1554_addr = 5'h8;
  assign tlb_entries_p1_v__T_1554_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1554_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1555_addr = 5'h9;
  assign tlb_entries_p1_v__T_1555_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1555_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1556_addr = 5'ha;
  assign tlb_entries_p1_v__T_1556_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1556_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1557_addr = 5'hb;
  assign tlb_entries_p1_v__T_1557_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1557_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1558_addr = 5'hc;
  assign tlb_entries_p1_v__T_1558_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1558_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1559_addr = 5'hd;
  assign tlb_entries_p1_v__T_1559_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1559_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1560_addr = 5'he;
  assign tlb_entries_p1_v__T_1560_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1560_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1561_addr = 5'hf;
  assign tlb_entries_p1_v__T_1561_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1561_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1562_addr = 5'h10;
  assign tlb_entries_p1_v__T_1562_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1562_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1563_addr = 5'h11;
  assign tlb_entries_p1_v__T_1563_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1563_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1564_addr = 5'h12;
  assign tlb_entries_p1_v__T_1564_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1564_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1565_addr = 5'h13;
  assign tlb_entries_p1_v__T_1565_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1565_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1566_addr = 5'h14;
  assign tlb_entries_p1_v__T_1566_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1566_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1567_addr = 5'h15;
  assign tlb_entries_p1_v__T_1567_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1567_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1568_addr = 5'h16;
  assign tlb_entries_p1_v__T_1568_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1568_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1569_addr = 5'h17;
  assign tlb_entries_p1_v__T_1569_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1569_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1570_addr = 5'h18;
  assign tlb_entries_p1_v__T_1570_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1570_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1571_addr = 5'h19;
  assign tlb_entries_p1_v__T_1571_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1571_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1572_addr = 5'h1a;
  assign tlb_entries_p1_v__T_1572_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1572_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1573_addr = 5'h1b;
  assign tlb_entries_p1_v__T_1573_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1573_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1574_addr = 5'h1c;
  assign tlb_entries_p1_v__T_1574_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1574_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1575_addr = 5'h1d;
  assign tlb_entries_p1_v__T_1575_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1575_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1576_addr = 5'h1e;
  assign tlb_entries_p1_v__T_1576_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1576_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v__T_1577_addr = 5'h1f;
  assign tlb_entries_p1_v__T_1577_data = tlb_entries_p1_v[tlb_entries_p1_v__T_1577_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_0_r_addr = 5'h0;
  assign tlb_entries_p1_v_tlb_entry_ports_0_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_0_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_1_r_addr = 5'h1;
  assign tlb_entries_p1_v_tlb_entry_ports_1_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_1_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_2_r_addr = 5'h2;
  assign tlb_entries_p1_v_tlb_entry_ports_2_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_2_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_3_r_addr = 5'h3;
  assign tlb_entries_p1_v_tlb_entry_ports_3_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_3_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_4_r_addr = 5'h4;
  assign tlb_entries_p1_v_tlb_entry_ports_4_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_4_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_5_r_addr = 5'h5;
  assign tlb_entries_p1_v_tlb_entry_ports_5_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_5_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_6_r_addr = 5'h6;
  assign tlb_entries_p1_v_tlb_entry_ports_6_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_6_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_7_r_addr = 5'h7;
  assign tlb_entries_p1_v_tlb_entry_ports_7_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_7_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_8_r_addr = 5'h8;
  assign tlb_entries_p1_v_tlb_entry_ports_8_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_8_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_9_r_addr = 5'h9;
  assign tlb_entries_p1_v_tlb_entry_ports_9_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_9_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_10_r_addr = 5'ha;
  assign tlb_entries_p1_v_tlb_entry_ports_10_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_10_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_11_r_addr = 5'hb;
  assign tlb_entries_p1_v_tlb_entry_ports_11_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_11_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_12_r_addr = 5'hc;
  assign tlb_entries_p1_v_tlb_entry_ports_12_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_12_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_13_r_addr = 5'hd;
  assign tlb_entries_p1_v_tlb_entry_ports_13_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_13_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_14_r_addr = 5'he;
  assign tlb_entries_p1_v_tlb_entry_ports_14_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_14_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_15_r_addr = 5'hf;
  assign tlb_entries_p1_v_tlb_entry_ports_15_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_15_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_16_r_addr = 5'h10;
  assign tlb_entries_p1_v_tlb_entry_ports_16_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_16_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_17_r_addr = 5'h11;
  assign tlb_entries_p1_v_tlb_entry_ports_17_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_17_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_18_r_addr = 5'h12;
  assign tlb_entries_p1_v_tlb_entry_ports_18_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_18_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_19_r_addr = 5'h13;
  assign tlb_entries_p1_v_tlb_entry_ports_19_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_19_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_20_r_addr = 5'h14;
  assign tlb_entries_p1_v_tlb_entry_ports_20_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_20_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_21_r_addr = 5'h15;
  assign tlb_entries_p1_v_tlb_entry_ports_21_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_21_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_22_r_addr = 5'h16;
  assign tlb_entries_p1_v_tlb_entry_ports_22_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_22_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_23_r_addr = 5'h17;
  assign tlb_entries_p1_v_tlb_entry_ports_23_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_23_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_24_r_addr = 5'h18;
  assign tlb_entries_p1_v_tlb_entry_ports_24_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_24_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_25_r_addr = 5'h19;
  assign tlb_entries_p1_v_tlb_entry_ports_25_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_25_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_26_r_addr = 5'h1a;
  assign tlb_entries_p1_v_tlb_entry_ports_26_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_26_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_27_r_addr = 5'h1b;
  assign tlb_entries_p1_v_tlb_entry_ports_27_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_27_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_28_r_addr = 5'h1c;
  assign tlb_entries_p1_v_tlb_entry_ports_28_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_28_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_29_r_addr = 5'h1d;
  assign tlb_entries_p1_v_tlb_entry_ports_29_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_29_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_30_r_addr = 5'h1e;
  assign tlb_entries_p1_v_tlb_entry_ports_30_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_30_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_31_r_addr = 5'h1f;
  assign tlb_entries_p1_v_tlb_entry_ports_31_r_data = tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_31_r_addr]; // @[tlb.scala 45:24]
  assign tlb_entries_p1_v_tlb_entry_ports_0_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_0_w_addr = 5'h0;
  assign tlb_entries_p1_v_tlb_entry_ports_0_w_mask = _T_3545 & _T_3546;
  assign tlb_entries_p1_v_tlb_entry_ports_0_w_en = _T_3545 & _T_3546;
  assign tlb_entries_p1_v_tlb_entry_ports_1_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_1_w_addr = 5'h1;
  assign tlb_entries_p1_v_tlb_entry_ports_1_w_mask = _T_3545 & _T_3547;
  assign tlb_entries_p1_v_tlb_entry_ports_1_w_en = _T_3545 & _T_3547;
  assign tlb_entries_p1_v_tlb_entry_ports_2_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_2_w_addr = 5'h2;
  assign tlb_entries_p1_v_tlb_entry_ports_2_w_mask = _T_3545 & _T_3548;
  assign tlb_entries_p1_v_tlb_entry_ports_2_w_en = _T_3545 & _T_3548;
  assign tlb_entries_p1_v_tlb_entry_ports_3_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_3_w_addr = 5'h3;
  assign tlb_entries_p1_v_tlb_entry_ports_3_w_mask = _T_3545 & _T_3549;
  assign tlb_entries_p1_v_tlb_entry_ports_3_w_en = _T_3545 & _T_3549;
  assign tlb_entries_p1_v_tlb_entry_ports_4_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_4_w_addr = 5'h4;
  assign tlb_entries_p1_v_tlb_entry_ports_4_w_mask = _T_3545 & _T_3550;
  assign tlb_entries_p1_v_tlb_entry_ports_4_w_en = _T_3545 & _T_3550;
  assign tlb_entries_p1_v_tlb_entry_ports_5_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_5_w_addr = 5'h5;
  assign tlb_entries_p1_v_tlb_entry_ports_5_w_mask = _T_3545 & _T_3551;
  assign tlb_entries_p1_v_tlb_entry_ports_5_w_en = _T_3545 & _T_3551;
  assign tlb_entries_p1_v_tlb_entry_ports_6_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_6_w_addr = 5'h6;
  assign tlb_entries_p1_v_tlb_entry_ports_6_w_mask = _T_3545 & _T_3552;
  assign tlb_entries_p1_v_tlb_entry_ports_6_w_en = _T_3545 & _T_3552;
  assign tlb_entries_p1_v_tlb_entry_ports_7_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_7_w_addr = 5'h7;
  assign tlb_entries_p1_v_tlb_entry_ports_7_w_mask = _T_3545 & _T_3553;
  assign tlb_entries_p1_v_tlb_entry_ports_7_w_en = _T_3545 & _T_3553;
  assign tlb_entries_p1_v_tlb_entry_ports_8_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_8_w_addr = 5'h8;
  assign tlb_entries_p1_v_tlb_entry_ports_8_w_mask = _T_3545 & _T_3554;
  assign tlb_entries_p1_v_tlb_entry_ports_8_w_en = _T_3545 & _T_3554;
  assign tlb_entries_p1_v_tlb_entry_ports_9_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_9_w_addr = 5'h9;
  assign tlb_entries_p1_v_tlb_entry_ports_9_w_mask = _T_3545 & _T_3555;
  assign tlb_entries_p1_v_tlb_entry_ports_9_w_en = _T_3545 & _T_3555;
  assign tlb_entries_p1_v_tlb_entry_ports_10_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_10_w_addr = 5'ha;
  assign tlb_entries_p1_v_tlb_entry_ports_10_w_mask = _T_3545 & _T_3556;
  assign tlb_entries_p1_v_tlb_entry_ports_10_w_en = _T_3545 & _T_3556;
  assign tlb_entries_p1_v_tlb_entry_ports_11_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_11_w_addr = 5'hb;
  assign tlb_entries_p1_v_tlb_entry_ports_11_w_mask = _T_3545 & _T_3557;
  assign tlb_entries_p1_v_tlb_entry_ports_11_w_en = _T_3545 & _T_3557;
  assign tlb_entries_p1_v_tlb_entry_ports_12_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_12_w_addr = 5'hc;
  assign tlb_entries_p1_v_tlb_entry_ports_12_w_mask = _T_3545 & _T_3558;
  assign tlb_entries_p1_v_tlb_entry_ports_12_w_en = _T_3545 & _T_3558;
  assign tlb_entries_p1_v_tlb_entry_ports_13_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_13_w_addr = 5'hd;
  assign tlb_entries_p1_v_tlb_entry_ports_13_w_mask = _T_3545 & _T_3559;
  assign tlb_entries_p1_v_tlb_entry_ports_13_w_en = _T_3545 & _T_3559;
  assign tlb_entries_p1_v_tlb_entry_ports_14_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_14_w_addr = 5'he;
  assign tlb_entries_p1_v_tlb_entry_ports_14_w_mask = _T_3545 & _T_3560;
  assign tlb_entries_p1_v_tlb_entry_ports_14_w_en = _T_3545 & _T_3560;
  assign tlb_entries_p1_v_tlb_entry_ports_15_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_15_w_addr = 5'hf;
  assign tlb_entries_p1_v_tlb_entry_ports_15_w_mask = _T_3545 & _T_3561;
  assign tlb_entries_p1_v_tlb_entry_ports_15_w_en = _T_3545 & _T_3561;
  assign tlb_entries_p1_v_tlb_entry_ports_16_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_16_w_addr = 5'h10;
  assign tlb_entries_p1_v_tlb_entry_ports_16_w_mask = _T_3545 & _T_3562;
  assign tlb_entries_p1_v_tlb_entry_ports_16_w_en = _T_3545 & _T_3562;
  assign tlb_entries_p1_v_tlb_entry_ports_17_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_17_w_addr = 5'h11;
  assign tlb_entries_p1_v_tlb_entry_ports_17_w_mask = _T_3545 & _T_3563;
  assign tlb_entries_p1_v_tlb_entry_ports_17_w_en = _T_3545 & _T_3563;
  assign tlb_entries_p1_v_tlb_entry_ports_18_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_18_w_addr = 5'h12;
  assign tlb_entries_p1_v_tlb_entry_ports_18_w_mask = _T_3545 & _T_3564;
  assign tlb_entries_p1_v_tlb_entry_ports_18_w_en = _T_3545 & _T_3564;
  assign tlb_entries_p1_v_tlb_entry_ports_19_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_19_w_addr = 5'h13;
  assign tlb_entries_p1_v_tlb_entry_ports_19_w_mask = _T_3545 & _T_3565;
  assign tlb_entries_p1_v_tlb_entry_ports_19_w_en = _T_3545 & _T_3565;
  assign tlb_entries_p1_v_tlb_entry_ports_20_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_20_w_addr = 5'h14;
  assign tlb_entries_p1_v_tlb_entry_ports_20_w_mask = _T_3545 & _T_3566;
  assign tlb_entries_p1_v_tlb_entry_ports_20_w_en = _T_3545 & _T_3566;
  assign tlb_entries_p1_v_tlb_entry_ports_21_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_21_w_addr = 5'h15;
  assign tlb_entries_p1_v_tlb_entry_ports_21_w_mask = _T_3545 & _T_3567;
  assign tlb_entries_p1_v_tlb_entry_ports_21_w_en = _T_3545 & _T_3567;
  assign tlb_entries_p1_v_tlb_entry_ports_22_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_22_w_addr = 5'h16;
  assign tlb_entries_p1_v_tlb_entry_ports_22_w_mask = _T_3545 & _T_3568;
  assign tlb_entries_p1_v_tlb_entry_ports_22_w_en = _T_3545 & _T_3568;
  assign tlb_entries_p1_v_tlb_entry_ports_23_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_23_w_addr = 5'h17;
  assign tlb_entries_p1_v_tlb_entry_ports_23_w_mask = _T_3545 & _T_3569;
  assign tlb_entries_p1_v_tlb_entry_ports_23_w_en = _T_3545 & _T_3569;
  assign tlb_entries_p1_v_tlb_entry_ports_24_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_24_w_addr = 5'h18;
  assign tlb_entries_p1_v_tlb_entry_ports_24_w_mask = _T_3545 & _T_3570;
  assign tlb_entries_p1_v_tlb_entry_ports_24_w_en = _T_3545 & _T_3570;
  assign tlb_entries_p1_v_tlb_entry_ports_25_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_25_w_addr = 5'h19;
  assign tlb_entries_p1_v_tlb_entry_ports_25_w_mask = _T_3545 & _T_3571;
  assign tlb_entries_p1_v_tlb_entry_ports_25_w_en = _T_3545 & _T_3571;
  assign tlb_entries_p1_v_tlb_entry_ports_26_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_26_w_addr = 5'h1a;
  assign tlb_entries_p1_v_tlb_entry_ports_26_w_mask = _T_3545 & _T_3572;
  assign tlb_entries_p1_v_tlb_entry_ports_26_w_en = _T_3545 & _T_3572;
  assign tlb_entries_p1_v_tlb_entry_ports_27_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_27_w_addr = 5'h1b;
  assign tlb_entries_p1_v_tlb_entry_ports_27_w_mask = _T_3545 & _T_3573;
  assign tlb_entries_p1_v_tlb_entry_ports_27_w_en = _T_3545 & _T_3573;
  assign tlb_entries_p1_v_tlb_entry_ports_28_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_28_w_addr = 5'h1c;
  assign tlb_entries_p1_v_tlb_entry_ports_28_w_mask = _T_3545 & _T_3574;
  assign tlb_entries_p1_v_tlb_entry_ports_28_w_en = _T_3545 & _T_3574;
  assign tlb_entries_p1_v_tlb_entry_ports_29_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_29_w_addr = 5'h1d;
  assign tlb_entries_p1_v_tlb_entry_ports_29_w_mask = _T_3545 & _T_3575;
  assign tlb_entries_p1_v_tlb_entry_ports_29_w_en = _T_3545 & _T_3575;
  assign tlb_entries_p1_v_tlb_entry_ports_30_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_30_w_addr = 5'h1e;
  assign tlb_entries_p1_v_tlb_entry_ports_30_w_mask = _T_3545 & _T_3576;
  assign tlb_entries_p1_v_tlb_entry_ports_30_w_en = _T_3545 & _T_3576;
  assign tlb_entries_p1_v_tlb_entry_ports_31_w_data = io_wport_bits_entry_p1_v;
  assign tlb_entries_p1_v_tlb_entry_ports_31_w_addr = 5'h1f;
  assign tlb_entries_p1_v_tlb_entry_ports_31_w_mask = _T_3545 & _T_3577;
  assign tlb_entries_p1_v_tlb_entry_ports_31_w_en = _T_3545 & _T_3577;
  assign io_iaddr_req_ready = io_iaddr_resp_ready | _T_1529; // @[tlb.scala 160:19]
  assign io_iaddr_resp_valid = _T_4; // @[tlb.scala 161:20]
  assign io_iaddr_resp_bits_paddr = _T_1494 | _T_1492; // @[tlb.scala 162:25]
  assign io_iaddr_resp_bits_is_cached = _T_3_vaddr[31:29] != 3'h5; // @[tlb.scala 163:29]
  assign io_iaddr_resp_bits_ex_et = _T_1523 ? 5'h6 : _T_1508; // @[tlb.scala 164:22]
  assign io_iaddr_resp_bits_ex_code = _T_1523 ? 5'h4 : _T_1473_ex_code; // @[tlb.scala 164:22]
  assign io_iaddr_resp_bits_ex_addr = _T_3_vaddr; // @[tlb.scala 164:22]
  assign io_iaddr_resp_bits_ex_asid = _T_1523 ? 8'h0 : _T_1473_ex_asid; // @[tlb.scala 164:22]
  assign io_daddr_req_ready = 1'h1; // @[tlb.scala 160:19]
  assign io_daddr_resp_bits_paddr = _T_3035 | _T_3033; // @[tlb.scala 162:25]
  assign io_daddr_resp_bits_ex_et = _T_3064 ? 5'h6 : _T_3049; // @[tlb.scala 164:22]
  assign io_daddr_resp_bits_ex_code = _T_3064 ? _T_3069 : _T_3014_ex_code; // @[tlb.scala 164:22]
  assign io_daddr_resp_bits_ex_addr = _T_1544_vaddr; // @[tlb.scala 164:22]
  assign io_daddr_resp_bits_ex_asid = _T_3064 ? 8'h0 : _T_3014_ex_asid; // @[tlb.scala 164:22]
  assign io_rport_entry_pagemask = _T_3529[101:86]; // @[tlb.scala 190:18]
  assign io_rport_entry_vpn = _T_3529[85:67]; // @[tlb.scala 190:18]
  assign io_rport_entry_g = _T_3529[66]; // @[tlb.scala 190:18]
  assign io_rport_entry_asid = _T_3529[65:58]; // @[tlb.scala 190:18]
  assign io_rport_entry_p0_pfn = _T_3529[57:34]; // @[tlb.scala 190:18]
  assign io_rport_entry_p0_c = _T_3529[33:31]; // @[tlb.scala 190:18]
  assign io_rport_entry_p0_d = _T_3529[30]; // @[tlb.scala 190:18]
  assign io_rport_entry_p0_v = _T_3529[29]; // @[tlb.scala 190:18]
  assign io_rport_entry_p1_pfn = _T_3529[28:5]; // @[tlb.scala 190:18]
  assign io_rport_entry_p1_c = _T_3529[4:2]; // @[tlb.scala 190:18]
  assign io_rport_entry_p1_d = _T_3529[1]; // @[tlb.scala 190:18]
  assign io_rport_entry_p1_v = _T_3529[0]; // @[tlb.scala 190:18]
  assign io_pport_index_p = ~_T_3945; // @[tlb.scala 203:20]
  assign io_pport_index_index = _T_4040 | _T_4010; // @[tlb.scala 204:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_pagemask[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_vpn[initvar] = _RAND_1[18:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_g[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_asid[initvar] = _RAND_3[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p0_pfn[initvar] = _RAND_4[23:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p0_c[initvar] = _RAND_5[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p0_d[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p0_v[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p1_pfn[initvar] = _RAND_8[23:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p1_c[initvar] = _RAND_9[2:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p1_d[initvar] = _RAND_10[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    tlb_entries_p1_v[initvar] = _RAND_11[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_3_vaddr = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_3_len = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_3_is_aligned = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_4 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1544_func = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1544_vaddr = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1544_len = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1544_is_aligned = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tlb_entries_pagemask_tlb_entry_ports_0_w_en & tlb_entries_pagemask_tlb_entry_ports_0_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_0_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_1_w_en & tlb_entries_pagemask_tlb_entry_ports_1_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_1_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_2_w_en & tlb_entries_pagemask_tlb_entry_ports_2_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_2_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_3_w_en & tlb_entries_pagemask_tlb_entry_ports_3_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_3_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_4_w_en & tlb_entries_pagemask_tlb_entry_ports_4_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_4_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_5_w_en & tlb_entries_pagemask_tlb_entry_ports_5_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_5_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_6_w_en & tlb_entries_pagemask_tlb_entry_ports_6_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_6_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_7_w_en & tlb_entries_pagemask_tlb_entry_ports_7_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_7_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_8_w_en & tlb_entries_pagemask_tlb_entry_ports_8_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_8_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_9_w_en & tlb_entries_pagemask_tlb_entry_ports_9_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_9_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_10_w_en & tlb_entries_pagemask_tlb_entry_ports_10_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_10_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_11_w_en & tlb_entries_pagemask_tlb_entry_ports_11_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_11_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_12_w_en & tlb_entries_pagemask_tlb_entry_ports_12_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_12_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_13_w_en & tlb_entries_pagemask_tlb_entry_ports_13_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_13_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_14_w_en & tlb_entries_pagemask_tlb_entry_ports_14_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_14_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_15_w_en & tlb_entries_pagemask_tlb_entry_ports_15_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_15_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_16_w_en & tlb_entries_pagemask_tlb_entry_ports_16_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_16_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_17_w_en & tlb_entries_pagemask_tlb_entry_ports_17_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_17_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_18_w_en & tlb_entries_pagemask_tlb_entry_ports_18_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_18_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_19_w_en & tlb_entries_pagemask_tlb_entry_ports_19_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_19_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_20_w_en & tlb_entries_pagemask_tlb_entry_ports_20_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_20_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_21_w_en & tlb_entries_pagemask_tlb_entry_ports_21_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_21_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_22_w_en & tlb_entries_pagemask_tlb_entry_ports_22_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_22_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_23_w_en & tlb_entries_pagemask_tlb_entry_ports_23_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_23_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_24_w_en & tlb_entries_pagemask_tlb_entry_ports_24_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_24_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_25_w_en & tlb_entries_pagemask_tlb_entry_ports_25_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_25_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_26_w_en & tlb_entries_pagemask_tlb_entry_ports_26_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_26_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_27_w_en & tlb_entries_pagemask_tlb_entry_ports_27_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_27_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_28_w_en & tlb_entries_pagemask_tlb_entry_ports_28_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_28_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_29_w_en & tlb_entries_pagemask_tlb_entry_ports_29_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_29_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_30_w_en & tlb_entries_pagemask_tlb_entry_ports_30_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_30_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_pagemask_tlb_entry_ports_31_w_en & tlb_entries_pagemask_tlb_entry_ports_31_w_mask) begin
      tlb_entries_pagemask[tlb_entries_pagemask_tlb_entry_ports_31_w_addr] <= tlb_entries_pagemask_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_0_w_en & tlb_entries_vpn_tlb_entry_ports_0_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_0_w_addr] <= tlb_entries_vpn_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_1_w_en & tlb_entries_vpn_tlb_entry_ports_1_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_1_w_addr] <= tlb_entries_vpn_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_2_w_en & tlb_entries_vpn_tlb_entry_ports_2_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_2_w_addr] <= tlb_entries_vpn_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_3_w_en & tlb_entries_vpn_tlb_entry_ports_3_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_3_w_addr] <= tlb_entries_vpn_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_4_w_en & tlb_entries_vpn_tlb_entry_ports_4_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_4_w_addr] <= tlb_entries_vpn_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_5_w_en & tlb_entries_vpn_tlb_entry_ports_5_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_5_w_addr] <= tlb_entries_vpn_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_6_w_en & tlb_entries_vpn_tlb_entry_ports_6_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_6_w_addr] <= tlb_entries_vpn_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_7_w_en & tlb_entries_vpn_tlb_entry_ports_7_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_7_w_addr] <= tlb_entries_vpn_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_8_w_en & tlb_entries_vpn_tlb_entry_ports_8_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_8_w_addr] <= tlb_entries_vpn_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_9_w_en & tlb_entries_vpn_tlb_entry_ports_9_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_9_w_addr] <= tlb_entries_vpn_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_10_w_en & tlb_entries_vpn_tlb_entry_ports_10_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_10_w_addr] <= tlb_entries_vpn_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_11_w_en & tlb_entries_vpn_tlb_entry_ports_11_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_11_w_addr] <= tlb_entries_vpn_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_12_w_en & tlb_entries_vpn_tlb_entry_ports_12_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_12_w_addr] <= tlb_entries_vpn_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_13_w_en & tlb_entries_vpn_tlb_entry_ports_13_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_13_w_addr] <= tlb_entries_vpn_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_14_w_en & tlb_entries_vpn_tlb_entry_ports_14_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_14_w_addr] <= tlb_entries_vpn_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_15_w_en & tlb_entries_vpn_tlb_entry_ports_15_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_15_w_addr] <= tlb_entries_vpn_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_16_w_en & tlb_entries_vpn_tlb_entry_ports_16_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_16_w_addr] <= tlb_entries_vpn_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_17_w_en & tlb_entries_vpn_tlb_entry_ports_17_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_17_w_addr] <= tlb_entries_vpn_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_18_w_en & tlb_entries_vpn_tlb_entry_ports_18_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_18_w_addr] <= tlb_entries_vpn_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_19_w_en & tlb_entries_vpn_tlb_entry_ports_19_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_19_w_addr] <= tlb_entries_vpn_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_20_w_en & tlb_entries_vpn_tlb_entry_ports_20_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_20_w_addr] <= tlb_entries_vpn_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_21_w_en & tlb_entries_vpn_tlb_entry_ports_21_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_21_w_addr] <= tlb_entries_vpn_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_22_w_en & tlb_entries_vpn_tlb_entry_ports_22_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_22_w_addr] <= tlb_entries_vpn_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_23_w_en & tlb_entries_vpn_tlb_entry_ports_23_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_23_w_addr] <= tlb_entries_vpn_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_24_w_en & tlb_entries_vpn_tlb_entry_ports_24_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_24_w_addr] <= tlb_entries_vpn_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_25_w_en & tlb_entries_vpn_tlb_entry_ports_25_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_25_w_addr] <= tlb_entries_vpn_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_26_w_en & tlb_entries_vpn_tlb_entry_ports_26_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_26_w_addr] <= tlb_entries_vpn_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_27_w_en & tlb_entries_vpn_tlb_entry_ports_27_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_27_w_addr] <= tlb_entries_vpn_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_28_w_en & tlb_entries_vpn_tlb_entry_ports_28_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_28_w_addr] <= tlb_entries_vpn_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_29_w_en & tlb_entries_vpn_tlb_entry_ports_29_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_29_w_addr] <= tlb_entries_vpn_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_30_w_en & tlb_entries_vpn_tlb_entry_ports_30_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_30_w_addr] <= tlb_entries_vpn_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_vpn_tlb_entry_ports_31_w_en & tlb_entries_vpn_tlb_entry_ports_31_w_mask) begin
      tlb_entries_vpn[tlb_entries_vpn_tlb_entry_ports_31_w_addr] <= tlb_entries_vpn_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_0_w_en & tlb_entries_g_tlb_entry_ports_0_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_0_w_addr] <= tlb_entries_g_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_1_w_en & tlb_entries_g_tlb_entry_ports_1_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_1_w_addr] <= tlb_entries_g_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_2_w_en & tlb_entries_g_tlb_entry_ports_2_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_2_w_addr] <= tlb_entries_g_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_3_w_en & tlb_entries_g_tlb_entry_ports_3_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_3_w_addr] <= tlb_entries_g_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_4_w_en & tlb_entries_g_tlb_entry_ports_4_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_4_w_addr] <= tlb_entries_g_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_5_w_en & tlb_entries_g_tlb_entry_ports_5_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_5_w_addr] <= tlb_entries_g_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_6_w_en & tlb_entries_g_tlb_entry_ports_6_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_6_w_addr] <= tlb_entries_g_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_7_w_en & tlb_entries_g_tlb_entry_ports_7_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_7_w_addr] <= tlb_entries_g_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_8_w_en & tlb_entries_g_tlb_entry_ports_8_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_8_w_addr] <= tlb_entries_g_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_9_w_en & tlb_entries_g_tlb_entry_ports_9_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_9_w_addr] <= tlb_entries_g_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_10_w_en & tlb_entries_g_tlb_entry_ports_10_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_10_w_addr] <= tlb_entries_g_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_11_w_en & tlb_entries_g_tlb_entry_ports_11_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_11_w_addr] <= tlb_entries_g_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_12_w_en & tlb_entries_g_tlb_entry_ports_12_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_12_w_addr] <= tlb_entries_g_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_13_w_en & tlb_entries_g_tlb_entry_ports_13_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_13_w_addr] <= tlb_entries_g_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_14_w_en & tlb_entries_g_tlb_entry_ports_14_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_14_w_addr] <= tlb_entries_g_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_15_w_en & tlb_entries_g_tlb_entry_ports_15_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_15_w_addr] <= tlb_entries_g_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_16_w_en & tlb_entries_g_tlb_entry_ports_16_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_16_w_addr] <= tlb_entries_g_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_17_w_en & tlb_entries_g_tlb_entry_ports_17_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_17_w_addr] <= tlb_entries_g_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_18_w_en & tlb_entries_g_tlb_entry_ports_18_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_18_w_addr] <= tlb_entries_g_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_19_w_en & tlb_entries_g_tlb_entry_ports_19_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_19_w_addr] <= tlb_entries_g_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_20_w_en & tlb_entries_g_tlb_entry_ports_20_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_20_w_addr] <= tlb_entries_g_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_21_w_en & tlb_entries_g_tlb_entry_ports_21_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_21_w_addr] <= tlb_entries_g_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_22_w_en & tlb_entries_g_tlb_entry_ports_22_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_22_w_addr] <= tlb_entries_g_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_23_w_en & tlb_entries_g_tlb_entry_ports_23_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_23_w_addr] <= tlb_entries_g_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_24_w_en & tlb_entries_g_tlb_entry_ports_24_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_24_w_addr] <= tlb_entries_g_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_25_w_en & tlb_entries_g_tlb_entry_ports_25_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_25_w_addr] <= tlb_entries_g_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_26_w_en & tlb_entries_g_tlb_entry_ports_26_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_26_w_addr] <= tlb_entries_g_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_27_w_en & tlb_entries_g_tlb_entry_ports_27_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_27_w_addr] <= tlb_entries_g_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_28_w_en & tlb_entries_g_tlb_entry_ports_28_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_28_w_addr] <= tlb_entries_g_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_29_w_en & tlb_entries_g_tlb_entry_ports_29_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_29_w_addr] <= tlb_entries_g_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_30_w_en & tlb_entries_g_tlb_entry_ports_30_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_30_w_addr] <= tlb_entries_g_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_g_tlb_entry_ports_31_w_en & tlb_entries_g_tlb_entry_ports_31_w_mask) begin
      tlb_entries_g[tlb_entries_g_tlb_entry_ports_31_w_addr] <= tlb_entries_g_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_0_w_en & tlb_entries_asid_tlb_entry_ports_0_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_0_w_addr] <= tlb_entries_asid_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_1_w_en & tlb_entries_asid_tlb_entry_ports_1_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_1_w_addr] <= tlb_entries_asid_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_2_w_en & tlb_entries_asid_tlb_entry_ports_2_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_2_w_addr] <= tlb_entries_asid_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_3_w_en & tlb_entries_asid_tlb_entry_ports_3_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_3_w_addr] <= tlb_entries_asid_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_4_w_en & tlb_entries_asid_tlb_entry_ports_4_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_4_w_addr] <= tlb_entries_asid_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_5_w_en & tlb_entries_asid_tlb_entry_ports_5_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_5_w_addr] <= tlb_entries_asid_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_6_w_en & tlb_entries_asid_tlb_entry_ports_6_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_6_w_addr] <= tlb_entries_asid_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_7_w_en & tlb_entries_asid_tlb_entry_ports_7_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_7_w_addr] <= tlb_entries_asid_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_8_w_en & tlb_entries_asid_tlb_entry_ports_8_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_8_w_addr] <= tlb_entries_asid_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_9_w_en & tlb_entries_asid_tlb_entry_ports_9_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_9_w_addr] <= tlb_entries_asid_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_10_w_en & tlb_entries_asid_tlb_entry_ports_10_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_10_w_addr] <= tlb_entries_asid_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_11_w_en & tlb_entries_asid_tlb_entry_ports_11_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_11_w_addr] <= tlb_entries_asid_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_12_w_en & tlb_entries_asid_tlb_entry_ports_12_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_12_w_addr] <= tlb_entries_asid_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_13_w_en & tlb_entries_asid_tlb_entry_ports_13_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_13_w_addr] <= tlb_entries_asid_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_14_w_en & tlb_entries_asid_tlb_entry_ports_14_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_14_w_addr] <= tlb_entries_asid_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_15_w_en & tlb_entries_asid_tlb_entry_ports_15_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_15_w_addr] <= tlb_entries_asid_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_16_w_en & tlb_entries_asid_tlb_entry_ports_16_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_16_w_addr] <= tlb_entries_asid_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_17_w_en & tlb_entries_asid_tlb_entry_ports_17_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_17_w_addr] <= tlb_entries_asid_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_18_w_en & tlb_entries_asid_tlb_entry_ports_18_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_18_w_addr] <= tlb_entries_asid_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_19_w_en & tlb_entries_asid_tlb_entry_ports_19_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_19_w_addr] <= tlb_entries_asid_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_20_w_en & tlb_entries_asid_tlb_entry_ports_20_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_20_w_addr] <= tlb_entries_asid_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_21_w_en & tlb_entries_asid_tlb_entry_ports_21_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_21_w_addr] <= tlb_entries_asid_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_22_w_en & tlb_entries_asid_tlb_entry_ports_22_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_22_w_addr] <= tlb_entries_asid_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_23_w_en & tlb_entries_asid_tlb_entry_ports_23_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_23_w_addr] <= tlb_entries_asid_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_24_w_en & tlb_entries_asid_tlb_entry_ports_24_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_24_w_addr] <= tlb_entries_asid_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_25_w_en & tlb_entries_asid_tlb_entry_ports_25_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_25_w_addr] <= tlb_entries_asid_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_26_w_en & tlb_entries_asid_tlb_entry_ports_26_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_26_w_addr] <= tlb_entries_asid_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_27_w_en & tlb_entries_asid_tlb_entry_ports_27_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_27_w_addr] <= tlb_entries_asid_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_28_w_en & tlb_entries_asid_tlb_entry_ports_28_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_28_w_addr] <= tlb_entries_asid_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_29_w_en & tlb_entries_asid_tlb_entry_ports_29_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_29_w_addr] <= tlb_entries_asid_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_30_w_en & tlb_entries_asid_tlb_entry_ports_30_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_30_w_addr] <= tlb_entries_asid_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_asid_tlb_entry_ports_31_w_en & tlb_entries_asid_tlb_entry_ports_31_w_mask) begin
      tlb_entries_asid[tlb_entries_asid_tlb_entry_ports_31_w_addr] <= tlb_entries_asid_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_0_w_en & tlb_entries_p0_pfn_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_0_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_1_w_en & tlb_entries_p0_pfn_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_1_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_2_w_en & tlb_entries_p0_pfn_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_2_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_3_w_en & tlb_entries_p0_pfn_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_3_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_4_w_en & tlb_entries_p0_pfn_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_4_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_5_w_en & tlb_entries_p0_pfn_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_5_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_6_w_en & tlb_entries_p0_pfn_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_6_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_7_w_en & tlb_entries_p0_pfn_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_7_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_8_w_en & tlb_entries_p0_pfn_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_8_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_9_w_en & tlb_entries_p0_pfn_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_9_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_10_w_en & tlb_entries_p0_pfn_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_10_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_11_w_en & tlb_entries_p0_pfn_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_11_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_12_w_en & tlb_entries_p0_pfn_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_12_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_13_w_en & tlb_entries_p0_pfn_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_13_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_14_w_en & tlb_entries_p0_pfn_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_14_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_15_w_en & tlb_entries_p0_pfn_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_15_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_16_w_en & tlb_entries_p0_pfn_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_16_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_17_w_en & tlb_entries_p0_pfn_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_17_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_18_w_en & tlb_entries_p0_pfn_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_18_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_19_w_en & tlb_entries_p0_pfn_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_19_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_20_w_en & tlb_entries_p0_pfn_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_20_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_21_w_en & tlb_entries_p0_pfn_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_21_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_22_w_en & tlb_entries_p0_pfn_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_22_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_23_w_en & tlb_entries_p0_pfn_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_23_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_24_w_en & tlb_entries_p0_pfn_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_24_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_25_w_en & tlb_entries_p0_pfn_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_25_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_26_w_en & tlb_entries_p0_pfn_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_26_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_27_w_en & tlb_entries_p0_pfn_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_27_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_28_w_en & tlb_entries_p0_pfn_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_28_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_29_w_en & tlb_entries_p0_pfn_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_29_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_30_w_en & tlb_entries_p0_pfn_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_30_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_pfn_tlb_entry_ports_31_w_en & tlb_entries_p0_pfn_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p0_pfn[tlb_entries_p0_pfn_tlb_entry_ports_31_w_addr] <= tlb_entries_p0_pfn_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_0_w_en & tlb_entries_p0_c_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_0_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_1_w_en & tlb_entries_p0_c_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_1_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_2_w_en & tlb_entries_p0_c_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_2_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_3_w_en & tlb_entries_p0_c_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_3_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_4_w_en & tlb_entries_p0_c_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_4_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_5_w_en & tlb_entries_p0_c_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_5_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_6_w_en & tlb_entries_p0_c_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_6_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_7_w_en & tlb_entries_p0_c_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_7_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_8_w_en & tlb_entries_p0_c_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_8_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_9_w_en & tlb_entries_p0_c_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_9_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_10_w_en & tlb_entries_p0_c_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_10_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_11_w_en & tlb_entries_p0_c_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_11_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_12_w_en & tlb_entries_p0_c_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_12_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_13_w_en & tlb_entries_p0_c_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_13_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_14_w_en & tlb_entries_p0_c_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_14_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_15_w_en & tlb_entries_p0_c_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_15_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_16_w_en & tlb_entries_p0_c_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_16_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_17_w_en & tlb_entries_p0_c_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_17_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_18_w_en & tlb_entries_p0_c_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_18_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_19_w_en & tlb_entries_p0_c_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_19_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_20_w_en & tlb_entries_p0_c_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_20_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_21_w_en & tlb_entries_p0_c_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_21_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_22_w_en & tlb_entries_p0_c_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_22_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_23_w_en & tlb_entries_p0_c_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_23_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_24_w_en & tlb_entries_p0_c_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_24_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_25_w_en & tlb_entries_p0_c_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_25_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_26_w_en & tlb_entries_p0_c_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_26_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_27_w_en & tlb_entries_p0_c_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_27_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_28_w_en & tlb_entries_p0_c_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_28_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_29_w_en & tlb_entries_p0_c_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_29_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_30_w_en & tlb_entries_p0_c_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_30_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_c_tlb_entry_ports_31_w_en & tlb_entries_p0_c_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p0_c[tlb_entries_p0_c_tlb_entry_ports_31_w_addr] <= tlb_entries_p0_c_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_0_w_en & tlb_entries_p0_d_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_0_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_1_w_en & tlb_entries_p0_d_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_1_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_2_w_en & tlb_entries_p0_d_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_2_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_3_w_en & tlb_entries_p0_d_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_3_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_4_w_en & tlb_entries_p0_d_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_4_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_5_w_en & tlb_entries_p0_d_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_5_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_6_w_en & tlb_entries_p0_d_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_6_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_7_w_en & tlb_entries_p0_d_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_7_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_8_w_en & tlb_entries_p0_d_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_8_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_9_w_en & tlb_entries_p0_d_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_9_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_10_w_en & tlb_entries_p0_d_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_10_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_11_w_en & tlb_entries_p0_d_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_11_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_12_w_en & tlb_entries_p0_d_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_12_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_13_w_en & tlb_entries_p0_d_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_13_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_14_w_en & tlb_entries_p0_d_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_14_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_15_w_en & tlb_entries_p0_d_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_15_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_16_w_en & tlb_entries_p0_d_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_16_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_17_w_en & tlb_entries_p0_d_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_17_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_18_w_en & tlb_entries_p0_d_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_18_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_19_w_en & tlb_entries_p0_d_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_19_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_20_w_en & tlb_entries_p0_d_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_20_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_21_w_en & tlb_entries_p0_d_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_21_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_22_w_en & tlb_entries_p0_d_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_22_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_23_w_en & tlb_entries_p0_d_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_23_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_24_w_en & tlb_entries_p0_d_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_24_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_25_w_en & tlb_entries_p0_d_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_25_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_26_w_en & tlb_entries_p0_d_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_26_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_27_w_en & tlb_entries_p0_d_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_27_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_28_w_en & tlb_entries_p0_d_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_28_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_29_w_en & tlb_entries_p0_d_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_29_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_30_w_en & tlb_entries_p0_d_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_30_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_d_tlb_entry_ports_31_w_en & tlb_entries_p0_d_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p0_d[tlb_entries_p0_d_tlb_entry_ports_31_w_addr] <= tlb_entries_p0_d_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_0_w_en & tlb_entries_p0_v_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_0_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_1_w_en & tlb_entries_p0_v_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_1_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_2_w_en & tlb_entries_p0_v_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_2_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_3_w_en & tlb_entries_p0_v_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_3_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_4_w_en & tlb_entries_p0_v_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_4_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_5_w_en & tlb_entries_p0_v_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_5_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_6_w_en & tlb_entries_p0_v_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_6_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_7_w_en & tlb_entries_p0_v_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_7_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_8_w_en & tlb_entries_p0_v_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_8_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_9_w_en & tlb_entries_p0_v_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_9_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_10_w_en & tlb_entries_p0_v_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_10_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_11_w_en & tlb_entries_p0_v_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_11_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_12_w_en & tlb_entries_p0_v_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_12_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_13_w_en & tlb_entries_p0_v_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_13_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_14_w_en & tlb_entries_p0_v_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_14_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_15_w_en & tlb_entries_p0_v_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_15_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_16_w_en & tlb_entries_p0_v_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_16_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_17_w_en & tlb_entries_p0_v_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_17_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_18_w_en & tlb_entries_p0_v_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_18_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_19_w_en & tlb_entries_p0_v_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_19_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_20_w_en & tlb_entries_p0_v_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_20_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_21_w_en & tlb_entries_p0_v_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_21_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_22_w_en & tlb_entries_p0_v_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_22_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_23_w_en & tlb_entries_p0_v_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_23_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_24_w_en & tlb_entries_p0_v_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_24_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_25_w_en & tlb_entries_p0_v_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_25_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_26_w_en & tlb_entries_p0_v_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_26_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_27_w_en & tlb_entries_p0_v_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_27_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_28_w_en & tlb_entries_p0_v_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_28_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_29_w_en & tlb_entries_p0_v_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_29_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_30_w_en & tlb_entries_p0_v_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_30_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p0_v_tlb_entry_ports_31_w_en & tlb_entries_p0_v_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p0_v[tlb_entries_p0_v_tlb_entry_ports_31_w_addr] <= tlb_entries_p0_v_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_0_w_en & tlb_entries_p1_pfn_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_0_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_1_w_en & tlb_entries_p1_pfn_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_1_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_2_w_en & tlb_entries_p1_pfn_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_2_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_3_w_en & tlb_entries_p1_pfn_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_3_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_4_w_en & tlb_entries_p1_pfn_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_4_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_5_w_en & tlb_entries_p1_pfn_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_5_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_6_w_en & tlb_entries_p1_pfn_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_6_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_7_w_en & tlb_entries_p1_pfn_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_7_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_8_w_en & tlb_entries_p1_pfn_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_8_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_9_w_en & tlb_entries_p1_pfn_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_9_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_10_w_en & tlb_entries_p1_pfn_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_10_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_11_w_en & tlb_entries_p1_pfn_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_11_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_12_w_en & tlb_entries_p1_pfn_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_12_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_13_w_en & tlb_entries_p1_pfn_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_13_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_14_w_en & tlb_entries_p1_pfn_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_14_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_15_w_en & tlb_entries_p1_pfn_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_15_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_16_w_en & tlb_entries_p1_pfn_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_16_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_17_w_en & tlb_entries_p1_pfn_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_17_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_18_w_en & tlb_entries_p1_pfn_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_18_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_19_w_en & tlb_entries_p1_pfn_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_19_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_20_w_en & tlb_entries_p1_pfn_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_20_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_21_w_en & tlb_entries_p1_pfn_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_21_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_22_w_en & tlb_entries_p1_pfn_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_22_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_23_w_en & tlb_entries_p1_pfn_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_23_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_24_w_en & tlb_entries_p1_pfn_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_24_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_25_w_en & tlb_entries_p1_pfn_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_25_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_26_w_en & tlb_entries_p1_pfn_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_26_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_27_w_en & tlb_entries_p1_pfn_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_27_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_28_w_en & tlb_entries_p1_pfn_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_28_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_29_w_en & tlb_entries_p1_pfn_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_29_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_30_w_en & tlb_entries_p1_pfn_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_30_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_pfn_tlb_entry_ports_31_w_en & tlb_entries_p1_pfn_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p1_pfn[tlb_entries_p1_pfn_tlb_entry_ports_31_w_addr] <= tlb_entries_p1_pfn_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_0_w_en & tlb_entries_p1_c_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_0_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_1_w_en & tlb_entries_p1_c_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_1_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_2_w_en & tlb_entries_p1_c_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_2_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_3_w_en & tlb_entries_p1_c_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_3_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_4_w_en & tlb_entries_p1_c_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_4_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_5_w_en & tlb_entries_p1_c_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_5_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_6_w_en & tlb_entries_p1_c_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_6_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_7_w_en & tlb_entries_p1_c_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_7_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_8_w_en & tlb_entries_p1_c_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_8_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_9_w_en & tlb_entries_p1_c_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_9_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_10_w_en & tlb_entries_p1_c_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_10_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_11_w_en & tlb_entries_p1_c_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_11_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_12_w_en & tlb_entries_p1_c_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_12_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_13_w_en & tlb_entries_p1_c_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_13_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_14_w_en & tlb_entries_p1_c_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_14_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_15_w_en & tlb_entries_p1_c_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_15_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_16_w_en & tlb_entries_p1_c_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_16_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_17_w_en & tlb_entries_p1_c_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_17_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_18_w_en & tlb_entries_p1_c_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_18_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_19_w_en & tlb_entries_p1_c_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_19_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_20_w_en & tlb_entries_p1_c_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_20_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_21_w_en & tlb_entries_p1_c_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_21_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_22_w_en & tlb_entries_p1_c_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_22_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_23_w_en & tlb_entries_p1_c_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_23_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_24_w_en & tlb_entries_p1_c_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_24_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_25_w_en & tlb_entries_p1_c_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_25_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_26_w_en & tlb_entries_p1_c_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_26_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_27_w_en & tlb_entries_p1_c_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_27_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_28_w_en & tlb_entries_p1_c_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_28_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_29_w_en & tlb_entries_p1_c_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_29_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_30_w_en & tlb_entries_p1_c_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_30_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_c_tlb_entry_ports_31_w_en & tlb_entries_p1_c_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p1_c[tlb_entries_p1_c_tlb_entry_ports_31_w_addr] <= tlb_entries_p1_c_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_0_w_en & tlb_entries_p1_d_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_0_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_1_w_en & tlb_entries_p1_d_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_1_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_2_w_en & tlb_entries_p1_d_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_2_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_3_w_en & tlb_entries_p1_d_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_3_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_4_w_en & tlb_entries_p1_d_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_4_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_5_w_en & tlb_entries_p1_d_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_5_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_6_w_en & tlb_entries_p1_d_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_6_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_7_w_en & tlb_entries_p1_d_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_7_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_8_w_en & tlb_entries_p1_d_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_8_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_9_w_en & tlb_entries_p1_d_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_9_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_10_w_en & tlb_entries_p1_d_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_10_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_11_w_en & tlb_entries_p1_d_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_11_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_12_w_en & tlb_entries_p1_d_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_12_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_13_w_en & tlb_entries_p1_d_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_13_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_14_w_en & tlb_entries_p1_d_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_14_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_15_w_en & tlb_entries_p1_d_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_15_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_16_w_en & tlb_entries_p1_d_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_16_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_17_w_en & tlb_entries_p1_d_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_17_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_18_w_en & tlb_entries_p1_d_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_18_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_19_w_en & tlb_entries_p1_d_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_19_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_20_w_en & tlb_entries_p1_d_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_20_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_21_w_en & tlb_entries_p1_d_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_21_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_22_w_en & tlb_entries_p1_d_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_22_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_23_w_en & tlb_entries_p1_d_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_23_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_24_w_en & tlb_entries_p1_d_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_24_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_25_w_en & tlb_entries_p1_d_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_25_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_26_w_en & tlb_entries_p1_d_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_26_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_27_w_en & tlb_entries_p1_d_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_27_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_28_w_en & tlb_entries_p1_d_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_28_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_29_w_en & tlb_entries_p1_d_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_29_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_30_w_en & tlb_entries_p1_d_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_30_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_d_tlb_entry_ports_31_w_en & tlb_entries_p1_d_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p1_d[tlb_entries_p1_d_tlb_entry_ports_31_w_addr] <= tlb_entries_p1_d_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_0_w_en & tlb_entries_p1_v_tlb_entry_ports_0_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_0_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_0_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_1_w_en & tlb_entries_p1_v_tlb_entry_ports_1_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_1_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_1_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_2_w_en & tlb_entries_p1_v_tlb_entry_ports_2_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_2_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_2_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_3_w_en & tlb_entries_p1_v_tlb_entry_ports_3_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_3_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_3_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_4_w_en & tlb_entries_p1_v_tlb_entry_ports_4_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_4_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_4_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_5_w_en & tlb_entries_p1_v_tlb_entry_ports_5_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_5_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_5_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_6_w_en & tlb_entries_p1_v_tlb_entry_ports_6_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_6_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_6_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_7_w_en & tlb_entries_p1_v_tlb_entry_ports_7_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_7_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_7_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_8_w_en & tlb_entries_p1_v_tlb_entry_ports_8_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_8_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_8_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_9_w_en & tlb_entries_p1_v_tlb_entry_ports_9_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_9_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_9_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_10_w_en & tlb_entries_p1_v_tlb_entry_ports_10_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_10_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_10_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_11_w_en & tlb_entries_p1_v_tlb_entry_ports_11_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_11_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_11_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_12_w_en & tlb_entries_p1_v_tlb_entry_ports_12_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_12_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_12_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_13_w_en & tlb_entries_p1_v_tlb_entry_ports_13_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_13_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_13_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_14_w_en & tlb_entries_p1_v_tlb_entry_ports_14_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_14_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_14_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_15_w_en & tlb_entries_p1_v_tlb_entry_ports_15_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_15_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_15_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_16_w_en & tlb_entries_p1_v_tlb_entry_ports_16_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_16_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_16_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_17_w_en & tlb_entries_p1_v_tlb_entry_ports_17_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_17_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_17_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_18_w_en & tlb_entries_p1_v_tlb_entry_ports_18_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_18_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_18_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_19_w_en & tlb_entries_p1_v_tlb_entry_ports_19_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_19_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_19_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_20_w_en & tlb_entries_p1_v_tlb_entry_ports_20_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_20_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_20_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_21_w_en & tlb_entries_p1_v_tlb_entry_ports_21_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_21_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_21_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_22_w_en & tlb_entries_p1_v_tlb_entry_ports_22_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_22_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_22_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_23_w_en & tlb_entries_p1_v_tlb_entry_ports_23_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_23_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_23_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_24_w_en & tlb_entries_p1_v_tlb_entry_ports_24_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_24_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_24_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_25_w_en & tlb_entries_p1_v_tlb_entry_ports_25_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_25_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_25_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_26_w_en & tlb_entries_p1_v_tlb_entry_ports_26_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_26_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_26_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_27_w_en & tlb_entries_p1_v_tlb_entry_ports_27_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_27_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_27_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_28_w_en & tlb_entries_p1_v_tlb_entry_ports_28_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_28_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_28_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_29_w_en & tlb_entries_p1_v_tlb_entry_ports_29_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_29_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_29_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_30_w_en & tlb_entries_p1_v_tlb_entry_ports_30_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_30_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_30_w_data; // @[tlb.scala 45:24]
    end
    if(tlb_entries_p1_v_tlb_entry_ports_31_w_en & tlb_entries_p1_v_tlb_entry_ports_31_w_mask) begin
      tlb_entries_p1_v[tlb_entries_p1_v_tlb_entry_ports_31_w_addr] <= tlb_entries_p1_v_tlb_entry_ports_31_w_data; // @[tlb.scala 45:24]
    end
    if (reset) begin
      _T_3_vaddr <= 32'h0;
    end else if (_T_1) begin
      _T_3_vaddr <= io_iaddr_req_bits_vaddr;
    end
    if (reset) begin
      _T_3_len <= 2'h0;
    end else if (_T_1) begin
      _T_3_len <= 2'h3;
    end
    if (reset) begin
      _T_3_is_aligned <= 1'h0;
    end else begin
      _T_3_is_aligned <= _GEN_0;
    end
    if (reset) begin
      _T_4 <= 1'h0;
    end else if (_T_1538) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= _GEN_196;
    end
    if (reset) begin
      _T_1544_func <= 1'h0;
    end else if (_T_1542) begin
      _T_1544_func <= io_daddr_req_bits_func;
    end
    if (reset) begin
      _T_1544_vaddr <= 32'h0;
    end else if (_T_1542) begin
      _T_1544_vaddr <= io_daddr_req_bits_vaddr;
    end
    if (reset) begin
      _T_1544_len <= 2'h0;
    end else if (_T_1542) begin
      _T_1544_len <= io_daddr_req_bits_len;
    end
    if (reset) begin
      _T_1544_is_aligned <= 1'h0;
    end else if (_T_1542) begin
      _T_1544_is_aligned <= io_daddr_req_bits_is_aligned;
    end
  end
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [7:0]  io_enq_bits_wb_id,
  input  [31:0] io_enq_bits_wb_pc,
  input  [5:0]  io_enq_bits_wb_instr_op,
  input  [4:0]  io_enq_bits_wb_instr_rs_idx,
  input  [4:0]  io_enq_bits_wb_instr_rt_idx,
  input  [4:0]  io_enq_bits_wb_instr_rd_idx,
  input  [4:0]  io_enq_bits_wb_instr_shamt,
  input  [5:0]  io_enq_bits_wb_instr_func,
  input  [4:0]  io_enq_bits_wb_rd_idx,
  input         io_enq_bits_wb_ip7,
  input         io_enq_bits_wb_is_br,
  input  [31:0] io_enq_bits_wb_npc,
  input  [4:0]  io_enq_bits_ops_fu_op,
  input  [31:0] io_enq_bits_ops_op1,
  input  [31:0] io_enq_bits_ops_op2,
  input         io_deq_ready,
  output        io_deq_valid,
  output [7:0]  io_deq_bits_wb_id,
  output [31:0] io_deq_bits_wb_pc,
  output [5:0]  io_deq_bits_wb_instr_op,
  output [4:0]  io_deq_bits_wb_instr_rs_idx,
  output [4:0]  io_deq_bits_wb_instr_rt_idx,
  output [4:0]  io_deq_bits_wb_instr_rd_idx,
  output [4:0]  io_deq_bits_wb_instr_shamt,
  output [5:0]  io_deq_bits_wb_instr_func,
  output [4:0]  io_deq_bits_wb_rd_idx,
  output        io_deq_bits_wb_ip7,
  output        io_deq_bits_wb_is_br,
  output [31:0] io_deq_bits_wb_npc,
  output [4:0]  io_deq_bits_ops_fu_op,
  output [31:0] io_deq_bits_ops_op1,
  output [31:0] io_deq_bits_ops_op2
);
  reg [7:0] _T_wb_id [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [7:0] _T_wb_id__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_id__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [7:0] _T_wb_id__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_id__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_id__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_id__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_wb_pc [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [31:0] _T_wb_pc__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_pc__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_3;
  wire [31:0] _T_wb_pc__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_pc__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_pc__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_pc__T_10_en; // @[Decoupled.scala 218:24]
  reg [5:0] _T_wb_instr_op [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_4;
  wire [5:0] _T_wb_instr_op__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_op__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_5;
  wire [5:0] _T_wb_instr_op__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_op__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_op__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_op__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_rs_idx [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_6;
  wire [4:0] _T_wb_instr_rs_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_rs_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_7;
  wire [4:0] _T_wb_instr_rs_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_rs_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rs_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rs_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_rt_idx [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_8;
  wire [4:0] _T_wb_instr_rt_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_rt_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_9;
  wire [4:0] _T_wb_instr_rt_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_rt_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rt_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rt_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_rd_idx [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_10;
  wire [4:0] _T_wb_instr_rd_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_rd_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_11;
  wire [4:0] _T_wb_instr_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_rd_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rd_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rd_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_shamt [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_12;
  wire [4:0] _T_wb_instr_shamt__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_shamt__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_13;
  wire [4:0] _T_wb_instr_shamt__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_shamt__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_shamt__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_shamt__T_10_en; // @[Decoupled.scala 218:24]
  reg [5:0] _T_wb_instr_func [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_14;
  wire [5:0] _T_wb_instr_func__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_func__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_15;
  wire [5:0] _T_wb_instr_func__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_instr_func__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_func__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_func__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_rd_idx [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_16;
  wire [4:0] _T_wb_rd_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_rd_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_17;
  wire [4:0] _T_wb_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_rd_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_rd_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_rd_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_wb_ip7 [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_18;
  wire  _T_wb_ip7__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_ip7__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_19;
  wire  _T_wb_ip7__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_ip7__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_ip7__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_ip7__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_wb_is_br [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_20;
  wire  _T_wb_is_br__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_is_br__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_21;
  wire  _T_wb_is_br__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_is_br__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_is_br__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_is_br__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_wb_npc [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_22;
  wire [31:0] _T_wb_npc__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_npc__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_23;
  wire [31:0] _T_wb_npc__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_wb_npc__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_npc__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_npc__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_ops_fu_op [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_24;
  wire [4:0] _T_ops_fu_op__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_ops_fu_op__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_25;
  wire [4:0] _T_ops_fu_op__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_ops_fu_op__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_ops_fu_op__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_ops_fu_op__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_ops_op1 [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_26;
  wire [31:0] _T_ops_op1__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_ops_op1__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_27;
  wire [31:0] _T_ops_op1__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_ops_op1__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_ops_op1__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_ops_op1__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_ops_op2 [0:2]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_28;
  wire [31:0] _T_ops_op2__T_18_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_ops_op2__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_29;
  wire [31:0] _T_ops_op2__T_10_data; // @[Decoupled.scala 218:24]
  wire [1:0] _T_ops_op2__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_ops_op2__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_ops_op2__T_10_en; // @[Decoupled.scala 218:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_30;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_31;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_32;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = value == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_12 = value + 2'h1; // @[Counter.scala 39:22]
  wire  wrap_1 = value_1 == 2'h2; // @[Counter.scala 38:24]
  wire [1:0] _T_14 = value_1 + 2'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_wb_id__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_id__T_18_data = _T_wb_id[_T_wb_id__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_id__T_18_data = _T_wb_id__T_18_addr >= 2'h3 ? _RAND_1[7:0] : _T_wb_id[_T_wb_id__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_id__T_10_data = io_enq_bits_wb_id;
  assign _T_wb_id__T_10_addr = value;
  assign _T_wb_id__T_10_mask = 1'h1;
  assign _T_wb_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_pc__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_pc__T_18_data = _T_wb_pc[_T_wb_pc__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_pc__T_18_data = _T_wb_pc__T_18_addr >= 2'h3 ? _RAND_3[31:0] : _T_wb_pc[_T_wb_pc__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_pc__T_10_data = io_enq_bits_wb_pc;
  assign _T_wb_pc__T_10_addr = value;
  assign _T_wb_pc__T_10_mask = 1'h1;
  assign _T_wb_pc__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_op__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_op__T_18_data = _T_wb_instr_op[_T_wb_instr_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_op__T_18_data = _T_wb_instr_op__T_18_addr >= 2'h3 ? _RAND_5[5:0] : _T_wb_instr_op[_T_wb_instr_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_op__T_10_data = io_enq_bits_wb_instr_op;
  assign _T_wb_instr_op__T_10_addr = value;
  assign _T_wb_instr_op__T_10_mask = 1'h1;
  assign _T_wb_instr_op__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_rs_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rs_idx__T_18_data = _T_wb_instr_rs_idx[_T_wb_instr_rs_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_rs_idx__T_18_data = _T_wb_instr_rs_idx__T_18_addr >= 2'h3 ? _RAND_7[4:0] : _T_wb_instr_rs_idx[_T_wb_instr_rs_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rs_idx__T_10_data = io_enq_bits_wb_instr_rs_idx;
  assign _T_wb_instr_rs_idx__T_10_addr = value;
  assign _T_wb_instr_rs_idx__T_10_mask = 1'h1;
  assign _T_wb_instr_rs_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_rt_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rt_idx__T_18_data = _T_wb_instr_rt_idx[_T_wb_instr_rt_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_rt_idx__T_18_data = _T_wb_instr_rt_idx__T_18_addr >= 2'h3 ? _RAND_9[4:0] : _T_wb_instr_rt_idx[_T_wb_instr_rt_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rt_idx__T_10_data = io_enq_bits_wb_instr_rt_idx;
  assign _T_wb_instr_rt_idx__T_10_addr = value;
  assign _T_wb_instr_rt_idx__T_10_mask = 1'h1;
  assign _T_wb_instr_rt_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_rd_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rd_idx__T_18_data = _T_wb_instr_rd_idx[_T_wb_instr_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_rd_idx__T_18_data = _T_wb_instr_rd_idx__T_18_addr >= 2'h3 ? _RAND_11[4:0] : _T_wb_instr_rd_idx[_T_wb_instr_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rd_idx__T_10_data = io_enq_bits_wb_instr_rd_idx;
  assign _T_wb_instr_rd_idx__T_10_addr = value;
  assign _T_wb_instr_rd_idx__T_10_mask = 1'h1;
  assign _T_wb_instr_rd_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_shamt__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_shamt__T_18_data = _T_wb_instr_shamt[_T_wb_instr_shamt__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_shamt__T_18_data = _T_wb_instr_shamt__T_18_addr >= 2'h3 ? _RAND_13[4:0] : _T_wb_instr_shamt[_T_wb_instr_shamt__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_shamt__T_10_data = io_enq_bits_wb_instr_shamt;
  assign _T_wb_instr_shamt__T_10_addr = value;
  assign _T_wb_instr_shamt__T_10_mask = 1'h1;
  assign _T_wb_instr_shamt__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_func__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_func__T_18_data = _T_wb_instr_func[_T_wb_instr_func__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_func__T_18_data = _T_wb_instr_func__T_18_addr >= 2'h3 ? _RAND_15[5:0] : _T_wb_instr_func[_T_wb_instr_func__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_func__T_10_data = io_enq_bits_wb_instr_func;
  assign _T_wb_instr_func__T_10_addr = value;
  assign _T_wb_instr_func__T_10_mask = 1'h1;
  assign _T_wb_instr_func__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_rd_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_rd_idx__T_18_data = _T_wb_rd_idx[_T_wb_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_rd_idx__T_18_data = _T_wb_rd_idx__T_18_addr >= 2'h3 ? _RAND_17[4:0] : _T_wb_rd_idx[_T_wb_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_rd_idx__T_10_data = io_enq_bits_wb_rd_idx;
  assign _T_wb_rd_idx__T_10_addr = value;
  assign _T_wb_rd_idx__T_10_mask = 1'h1;
  assign _T_wb_rd_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_ip7__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_ip7__T_18_data = _T_wb_ip7[_T_wb_ip7__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_ip7__T_18_data = _T_wb_ip7__T_18_addr >= 2'h3 ? _RAND_19[0:0] : _T_wb_ip7[_T_wb_ip7__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_ip7__T_10_data = io_enq_bits_wb_ip7;
  assign _T_wb_ip7__T_10_addr = value;
  assign _T_wb_ip7__T_10_mask = 1'h1;
  assign _T_wb_ip7__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_is_br__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_is_br__T_18_data = _T_wb_is_br[_T_wb_is_br__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_is_br__T_18_data = _T_wb_is_br__T_18_addr >= 2'h3 ? _RAND_21[0:0] : _T_wb_is_br[_T_wb_is_br__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_is_br__T_10_data = io_enq_bits_wb_is_br;
  assign _T_wb_is_br__T_10_addr = value;
  assign _T_wb_is_br__T_10_mask = 1'h1;
  assign _T_wb_is_br__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_npc__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_npc__T_18_data = _T_wb_npc[_T_wb_npc__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_npc__T_18_data = _T_wb_npc__T_18_addr >= 2'h3 ? _RAND_23[31:0] : _T_wb_npc[_T_wb_npc__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_npc__T_10_data = io_enq_bits_wb_npc;
  assign _T_wb_npc__T_10_addr = value;
  assign _T_wb_npc__T_10_mask = 1'h1;
  assign _T_wb_npc__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_ops_fu_op__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_ops_fu_op__T_18_data = _T_ops_fu_op[_T_ops_fu_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_ops_fu_op__T_18_data = _T_ops_fu_op__T_18_addr >= 2'h3 ? _RAND_25[4:0] : _T_ops_fu_op[_T_ops_fu_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_ops_fu_op__T_10_data = io_enq_bits_ops_fu_op;
  assign _T_ops_fu_op__T_10_addr = value;
  assign _T_ops_fu_op__T_10_mask = 1'h1;
  assign _T_ops_fu_op__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_ops_op1__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_ops_op1__T_18_data = _T_ops_op1[_T_ops_op1__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_ops_op1__T_18_data = _T_ops_op1__T_18_addr >= 2'h3 ? _RAND_27[31:0] : _T_ops_op1[_T_ops_op1__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_ops_op1__T_10_data = io_enq_bits_ops_op1;
  assign _T_ops_op1__T_10_addr = value;
  assign _T_ops_op1__T_10_mask = 1'h1;
  assign _T_ops_op1__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_ops_op2__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_ops_op2__T_18_data = _T_ops_op2[_T_ops_op2__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_ops_op2__T_18_data = _T_ops_op2__T_18_addr >= 2'h3 ? _RAND_29[31:0] : _T_ops_op2[_T_ops_op2__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_ops_op2__T_10_data = io_enq_bits_ops_op2;
  assign _T_ops_op2__T_10_addr = value;
  assign _T_ops_op2__T_10_mask = 1'h1;
  assign _T_ops_op2__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_wb_id = _T_wb_id__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_pc = _T_wb_pc__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_op = _T_wb_instr_op__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_rs_idx = _T_wb_instr_rs_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_rt_idx = _T_wb_instr_rt_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_rd_idx = _T_wb_instr_rd_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_shamt = _T_wb_instr_shamt__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_func = _T_wb_instr_func__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_rd_idx = _T_wb_rd_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_ip7 = _T_wb_ip7__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_is_br = _T_wb_is_br__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_npc = _T_wb_npc__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ops_fu_op = _T_ops_fu_op__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ops_op1 = _T_ops_op1__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ops_op2 = _T_ops_op2__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_id[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_pc[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_instr_op[initvar] = _RAND_4[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_instr_rs_idx[initvar] = _RAND_6[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_instr_rt_idx[initvar] = _RAND_8[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_instr_rd_idx[initvar] = _RAND_10[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_instr_shamt[initvar] = _RAND_12[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_instr_func[initvar] = _RAND_14[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_rd_idx[initvar] = _RAND_16[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_ip7[initvar] = _RAND_18[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {1{`RANDOM}};
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_is_br[initvar] = _RAND_20[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_wb_npc[initvar] = _RAND_22[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_23 = {1{`RANDOM}};
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_ops_fu_op[initvar] = _RAND_24[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  _RAND_26 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_ops_op1[initvar] = _RAND_26[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_27 = {1{`RANDOM}};
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_ops_op2[initvar] = _RAND_28[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  value = _RAND_30[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  value_1 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_wb_id__T_10_en & _T_wb_id__T_10_mask) begin
      _T_wb_id[_T_wb_id__T_10_addr] <= _T_wb_id__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_pc__T_10_en & _T_wb_pc__T_10_mask) begin
      _T_wb_pc[_T_wb_pc__T_10_addr] <= _T_wb_pc__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_op__T_10_en & _T_wb_instr_op__T_10_mask) begin
      _T_wb_instr_op[_T_wb_instr_op__T_10_addr] <= _T_wb_instr_op__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_rs_idx__T_10_en & _T_wb_instr_rs_idx__T_10_mask) begin
      _T_wb_instr_rs_idx[_T_wb_instr_rs_idx__T_10_addr] <= _T_wb_instr_rs_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_rt_idx__T_10_en & _T_wb_instr_rt_idx__T_10_mask) begin
      _T_wb_instr_rt_idx[_T_wb_instr_rt_idx__T_10_addr] <= _T_wb_instr_rt_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_rd_idx__T_10_en & _T_wb_instr_rd_idx__T_10_mask) begin
      _T_wb_instr_rd_idx[_T_wb_instr_rd_idx__T_10_addr] <= _T_wb_instr_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_shamt__T_10_en & _T_wb_instr_shamt__T_10_mask) begin
      _T_wb_instr_shamt[_T_wb_instr_shamt__T_10_addr] <= _T_wb_instr_shamt__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_func__T_10_en & _T_wb_instr_func__T_10_mask) begin
      _T_wb_instr_func[_T_wb_instr_func__T_10_addr] <= _T_wb_instr_func__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_rd_idx__T_10_en & _T_wb_rd_idx__T_10_mask) begin
      _T_wb_rd_idx[_T_wb_rd_idx__T_10_addr] <= _T_wb_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_ip7__T_10_en & _T_wb_ip7__T_10_mask) begin
      _T_wb_ip7[_T_wb_ip7__T_10_addr] <= _T_wb_ip7__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_is_br__T_10_en & _T_wb_is_br__T_10_mask) begin
      _T_wb_is_br[_T_wb_is_br__T_10_addr] <= _T_wb_is_br__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_npc__T_10_en & _T_wb_npc__T_10_mask) begin
      _T_wb_npc[_T_wb_npc__T_10_addr] <= _T_wb_npc__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_ops_fu_op__T_10_en & _T_ops_fu_op__T_10_mask) begin
      _T_ops_fu_op[_T_ops_fu_op__T_10_addr] <= _T_ops_fu_op__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_ops_op1__T_10_en & _T_ops_op1__T_10_mask) begin
      _T_ops_op1[_T_ops_op1__T_10_addr] <= _T_ops_op1__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_ops_op2__T_10_en & _T_ops_op2__T_10_mask) begin
      _T_ops_op2[_T_ops_op2__T_10_addr] <= _T_ops_op2__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (_T_6) begin
      if (wrap) begin
        value <= 2'h0;
      end else begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (_T_8) begin
      if (wrap_1) begin
        value_1 <= 2'h0;
      end else begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module LSU(
  input         clock,
  input         reset,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output        io_dmem_req_bits_is_cached,
  output [31:0] io_dmem_req_bits_addr,
  output [1:0]  io_dmem_req_bits_len,
  output [3:0]  io_dmem_req_bits_strb,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_func,
  output        io_dmem_resp_ready,
  input         io_dmem_resp_valid,
  input  [31:0] io_dmem_resp_bits_data,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_ip7,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  input  [4:0]  io_fu_in_bits_ops_fu_op,
  input  [31:0] io_fu_in_bits_ops_op1,
  input  [31:0] io_fu_in_bits_ops_op2,
  input         io_fu_in_bits_is_cached,
  output        io_fu_out_valid,
  output        io_fu_out_bits_v,
  output [7:0]  io_fu_out_bits_id,
  output [31:0] io_fu_out_bits_pc,
  output [5:0]  io_fu_out_bits_instr_op,
  output [4:0]  io_fu_out_bits_instr_rs_idx,
  output [4:0]  io_fu_out_bits_instr_rt_idx,
  output [4:0]  io_fu_out_bits_instr_rd_idx,
  output [4:0]  io_fu_out_bits_instr_shamt,
  output [5:0]  io_fu_out_bits_instr_func,
  output [4:0]  io_fu_out_bits_rd_idx,
  output        io_fu_out_bits_wen,
  output [31:0] io_fu_out_bits_data,
  output        io_fu_out_bits_ip7,
  output        io_fu_out_bits_is_br,
  output [31:0] io_fu_out_bits_npc,
  output        io_working
);
  wire  s2_datas_clock; // @[lsu.scala 95:24]
  wire  s2_datas_reset; // @[lsu.scala 95:24]
  wire  s2_datas_io_enq_ready; // @[lsu.scala 95:24]
  wire  s2_datas_io_enq_valid; // @[lsu.scala 95:24]
  wire [7:0] s2_datas_io_enq_bits_wb_id; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_enq_bits_wb_pc; // @[lsu.scala 95:24]
  wire [5:0] s2_datas_io_enq_bits_wb_instr_op; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_enq_bits_wb_instr_rs_idx; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_enq_bits_wb_instr_rt_idx; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_enq_bits_wb_instr_rd_idx; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_enq_bits_wb_instr_shamt; // @[lsu.scala 95:24]
  wire [5:0] s2_datas_io_enq_bits_wb_instr_func; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_enq_bits_wb_rd_idx; // @[lsu.scala 95:24]
  wire  s2_datas_io_enq_bits_wb_ip7; // @[lsu.scala 95:24]
  wire  s2_datas_io_enq_bits_wb_is_br; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_enq_bits_wb_npc; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_enq_bits_ops_fu_op; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_enq_bits_ops_op1; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_enq_bits_ops_op2; // @[lsu.scala 95:24]
  wire  s2_datas_io_deq_ready; // @[lsu.scala 95:24]
  wire  s2_datas_io_deq_valid; // @[lsu.scala 95:24]
  wire [7:0] s2_datas_io_deq_bits_wb_id; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_deq_bits_wb_pc; // @[lsu.scala 95:24]
  wire [5:0] s2_datas_io_deq_bits_wb_instr_op; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_deq_bits_wb_instr_rs_idx; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_deq_bits_wb_instr_rt_idx; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_deq_bits_wb_instr_rd_idx; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_deq_bits_wb_instr_shamt; // @[lsu.scala 95:24]
  wire [5:0] s2_datas_io_deq_bits_wb_instr_func; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_deq_bits_wb_rd_idx; // @[lsu.scala 95:24]
  wire  s2_datas_io_deq_bits_wb_ip7; // @[lsu.scala 95:24]
  wire  s2_datas_io_deq_bits_wb_is_br; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_deq_bits_wb_npc; // @[lsu.scala 95:24]
  wire [4:0] s2_datas_io_deq_bits_ops_fu_op; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_deq_bits_ops_op1; // @[lsu.scala 95:24]
  wire [31:0] s2_datas_io_deq_bits_ops_op2; // @[lsu.scala 95:24]
  wire  _T_30 = ~io_fu_in_valid; // @[lsu.scala 90:21]
  wire  s2_in_op_ext = io_fu_in_bits_ops_fu_op[0]; // @[lsu.scala 94:42]
  wire [1:0] s2_in_op_len = io_fu_in_bits_ops_fu_op[2:1]; // @[lsu.scala 94:42]
  wire  s2_in_op_align = io_fu_in_bits_ops_fu_op[4]; // @[lsu.scala 94:42]
  wire  _T_42 = ~s2_in_op_align; // @[lsu.scala 67:9]
  wire  _T_88 = ~s2_in_op_ext; // @[lsu.scala 67:23]
  wire  _T_89 = _T_42 & _T_88; // @[lsu.scala 67:16]
  wire [1:0] _T_90 = ~io_fu_in_bits_ops_op1[1:0]; // @[lsu.scala 68:18]
  wire [4:0] _T_91 = {_T_90, 3'h0}; // @[lsu.scala 68:23]
  wire [31:0] _T_92 = io_fu_in_bits_ops_op2 >> _T_91; // @[lsu.scala 68:14]
  wire [4:0] _T_93 = {io_fu_in_bits_ops_op1[1:0], 3'h0}; // @[lsu.scala 68:43]
  wire [62:0] _GEN_0 = {{31'd0}, io_fu_in_bits_ops_op2}; // @[lsu.scala 68:35]
  wire [62:0] _T_94 = _GEN_0 << _T_93; // @[lsu.scala 68:35]
  wire [62:0] _T_95 = _T_89 ? {{31'd0}, _T_92} : _T_94; // @[lsu.scala 67:8]
  wire [1:0] _T_96 = ~s2_in_op_len; // @[lsu.scala 44:23]
  wire [3:0] _T_97 = 4'hf >> _T_96; // @[lsu.scala 44:19]
  wire [6:0] _GEN_1 = {{3'd0}, _T_97}; // @[lsu.scala 44:30]
  wire [6:0] _T_99 = _GEN_1 << io_fu_in_bits_ops_op1[1:0]; // @[lsu.scala 44:30]
  wire [3:0] _T_103 = 4'hf >> _T_90; // @[lsu.scala 46:20]
  wire [6:0] _T_106 = 7'h78 >> _T_90; // @[lsu.scala 47:20]
  wire [6:0] _T_107 = _T_88 ? {{3'd0}, _T_103} : _T_106; // @[lsu.scala 45:8]
  wire [6:0] _T_108 = s2_in_op_align ? _T_99 : _T_107; // @[lsu.scala 43:30]
  wire [4:0] _T_110 = s2_datas_io_deq_bits_ops_fu_op;
  wire  s3_in_op_ext = _T_110[0]; // @[lsu.scala 112:42]
  wire [1:0] s3_in_op_len = _T_110[2:1]; // @[lsu.scala 112:42]
  wire  s3_in_op_func = _T_110[3]; // @[lsu.scala 112:42]
  wire  s3_in_op_align = _T_110[4]; // @[lsu.scala 112:42]
  wire [31:0] _T_115 = s3_in_op_align ? 32'h0 : s2_datas_io_deq_bits_ops_op2; // @[lsu.scala 114:32]
  wire [1:0] _T_117 = ~s3_in_op_len; // @[lsu.scala 44:23]
  wire [3:0] _T_118 = 4'hf >> _T_117; // @[lsu.scala 44:19]
  wire [6:0] _GEN_2 = {{3'd0}, _T_118}; // @[lsu.scala 44:30]
  wire [6:0] _T_120 = _GEN_2 << s2_datas_io_deq_bits_ops_op1[1:0]; // @[lsu.scala 44:30]
  wire  _T_121 = ~s3_in_op_ext; // @[lsu.scala 45:13]
  wire [1:0] _T_123 = ~s2_datas_io_deq_bits_ops_op1[1:0]; // @[lsu.scala 46:24]
  wire [3:0] _T_124 = 4'hf >> _T_123; // @[lsu.scala 46:20]
  wire [6:0] _T_127 = 7'h78 >> _T_123; // @[lsu.scala 47:20]
  wire [6:0] _T_128 = _T_121 ? {{3'd0}, _T_124} : _T_127; // @[lsu.scala 45:8]
  wire [6:0] _T_129 = s3_in_op_align ? _T_120 : _T_128; // @[lsu.scala 43:30]
  wire  _T_133 = _T_129[0]; // @[lsu.scala 50:60]
  wire  _T_136 = _T_129[1]; // @[lsu.scala 50:60]
  wire  _T_139 = _T_129[2]; // @[lsu.scala 50:60]
  wire  _T_142 = _T_129[3]; // @[lsu.scala 50:60]
  wire [7:0] _T_143 = {8{_T_142}}; // @[Cat.scala 29:58]
  wire [7:0] _T_144 = {8{_T_139}}; // @[Cat.scala 29:58]
  wire [7:0] _T_146 = {8{_T_136}}; // @[Cat.scala 29:58]
  wire [7:0] _T_147 = {8{_T_133}}; // @[Cat.scala 29:58]
  wire [31:0] _T_149 = {_T_147,_T_146,_T_144,_T_143}; // @[Cat.scala 29:58]
  wire [31:0] _T_153 = {{16'd0}, _T_149[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_155 = {_T_149[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_157 = _T_155 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_158 = _T_153 | _T_157; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{8'd0}, _T_158[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_163 = _GEN_3 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_165 = {_T_158[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_167 = _T_165 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_168 = _T_163 | _T_167; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_4 = {{4'd0}, _T_168[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_173 = _GEN_4 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_175 = {_T_168[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_177 = _T_175 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_178 = _T_173 | _T_177; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_5 = {{2'd0}, _T_178[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_183 = _GEN_5 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_185 = {_T_178[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_187 = _T_185 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_188 = _T_183 | _T_187; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_6 = {{1'd0}, _T_188[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_193 = _GEN_6 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_195 = {_T_188[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_197 = _T_195 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_198 = _T_193 | _T_197; // @[Bitwise.scala 103:39]
  wire  _T_199 = ~s3_in_op_align; // @[lsu.scala 55:21]
  wire  _T_201 = _T_199 & _T_121; // @[lsu.scala 55:28]
  wire [4:0] _T_203 = {_T_123, 3'h0}; // @[lsu.scala 56:23]
  wire [62:0] _GEN_7 = {{31'd0}, io_dmem_resp_bits_data}; // @[lsu.scala 56:12]
  wire [62:0] _T_204 = _GEN_7 << _T_203; // @[lsu.scala 56:12]
  wire [4:0] _T_205 = {s2_datas_io_deq_bits_ops_op1[1:0], 3'h0}; // @[lsu.scala 56:43]
  wire [31:0] _T_206 = io_dmem_resp_bits_data >> _T_205; // @[lsu.scala 56:35]
  wire [62:0] _T_207 = _T_201 ? _T_204 : {{31'd0}, _T_206}; // @[lsu.scala 55:20]
  wire [62:0] _GEN_8 = {{31'd0}, _T_198}; // @[lsu.scala 58:12]
  wire [62:0] _T_213 = _GEN_8 << _T_203; // @[lsu.scala 58:12]
  wire [31:0] _T_215 = _T_198 >> _T_205; // @[lsu.scala 58:35]
  wire [62:0] _T_216 = _T_201 ? _T_213 : {{31'd0}, _T_215}; // @[lsu.scala 57:20]
  wire [62:0] _T_217 = _T_207 & _T_216; // @[lsu.scala 63:12]
  wire [62:0] _T_218 = ~_T_216; // @[lsu.scala 63:32]
  wire [62:0] _GEN_9 = {{31'd0}, _T_115}; // @[lsu.scala 63:30]
  wire [62:0] _T_219 = _GEN_9 & _T_218; // @[lsu.scala 63:30]
  wire [62:0] ret_data = _T_217 | _T_219; // @[lsu.scala 63:21]
  wire  _T_220 = ~s3_in_op_func; // @[lsu.scala 118:37]
  wire [4:0] _T_223 = {s3_in_op_align,s3_in_op_func,s3_in_op_len,s3_in_op_ext}; // @[lsu.scala 118:59]
  wire  _T_224 = _T_223 == 5'h1f; // @[lsu.scala 118:66]
  wire  _T_239 = _T_223 == 5'h10; // @[lsu.scala 130:22]
  wire [7:0] _T_242 = ret_data[7:0]; // @[lsu.scala 130:60]
  wire [31:0] _T_243 = {{24{_T_242[7]}},_T_242}; // @[lsu.scala 130:73]
  wire  _T_247 = _T_223 == 5'h12; // @[lsu.scala 131:22]
  wire [15:0] _T_250 = ret_data[15:0]; // @[lsu.scala 131:61]
  wire [31:0] _T_251 = {{16{_T_250[15]}},_T_250}; // @[lsu.scala 131:74]
  wire [62:0] _T_252 = _T_247 ? {{31'd0}, _T_251} : ret_data; // @[Mux.scala 87:16]
  wire [62:0] _T_253 = _T_239 ? {{31'd0}, _T_243} : _T_252; // @[Mux.scala 87:16]
  wire [62:0] _T_254 = _T_224 ? 63'h1 : _T_253; // @[Mux.scala 87:16]
  Queue s2_datas ( // @[lsu.scala 95:24]
    .clock(s2_datas_clock),
    .reset(s2_datas_reset),
    .io_enq_ready(s2_datas_io_enq_ready),
    .io_enq_valid(s2_datas_io_enq_valid),
    .io_enq_bits_wb_id(s2_datas_io_enq_bits_wb_id),
    .io_enq_bits_wb_pc(s2_datas_io_enq_bits_wb_pc),
    .io_enq_bits_wb_instr_op(s2_datas_io_enq_bits_wb_instr_op),
    .io_enq_bits_wb_instr_rs_idx(s2_datas_io_enq_bits_wb_instr_rs_idx),
    .io_enq_bits_wb_instr_rt_idx(s2_datas_io_enq_bits_wb_instr_rt_idx),
    .io_enq_bits_wb_instr_rd_idx(s2_datas_io_enq_bits_wb_instr_rd_idx),
    .io_enq_bits_wb_instr_shamt(s2_datas_io_enq_bits_wb_instr_shamt),
    .io_enq_bits_wb_instr_func(s2_datas_io_enq_bits_wb_instr_func),
    .io_enq_bits_wb_rd_idx(s2_datas_io_enq_bits_wb_rd_idx),
    .io_enq_bits_wb_ip7(s2_datas_io_enq_bits_wb_ip7),
    .io_enq_bits_wb_is_br(s2_datas_io_enq_bits_wb_is_br),
    .io_enq_bits_wb_npc(s2_datas_io_enq_bits_wb_npc),
    .io_enq_bits_ops_fu_op(s2_datas_io_enq_bits_ops_fu_op),
    .io_enq_bits_ops_op1(s2_datas_io_enq_bits_ops_op1),
    .io_enq_bits_ops_op2(s2_datas_io_enq_bits_ops_op2),
    .io_deq_ready(s2_datas_io_deq_ready),
    .io_deq_valid(s2_datas_io_deq_valid),
    .io_deq_bits_wb_id(s2_datas_io_deq_bits_wb_id),
    .io_deq_bits_wb_pc(s2_datas_io_deq_bits_wb_pc),
    .io_deq_bits_wb_instr_op(s2_datas_io_deq_bits_wb_instr_op),
    .io_deq_bits_wb_instr_rs_idx(s2_datas_io_deq_bits_wb_instr_rs_idx),
    .io_deq_bits_wb_instr_rt_idx(s2_datas_io_deq_bits_wb_instr_rt_idx),
    .io_deq_bits_wb_instr_rd_idx(s2_datas_io_deq_bits_wb_instr_rd_idx),
    .io_deq_bits_wb_instr_shamt(s2_datas_io_deq_bits_wb_instr_shamt),
    .io_deq_bits_wb_instr_func(s2_datas_io_deq_bits_wb_instr_func),
    .io_deq_bits_wb_rd_idx(s2_datas_io_deq_bits_wb_rd_idx),
    .io_deq_bits_wb_ip7(s2_datas_io_deq_bits_wb_ip7),
    .io_deq_bits_wb_is_br(s2_datas_io_deq_bits_wb_is_br),
    .io_deq_bits_wb_npc(s2_datas_io_deq_bits_wb_npc),
    .io_deq_bits_ops_fu_op(s2_datas_io_deq_bits_ops_fu_op),
    .io_deq_bits_ops_op1(s2_datas_io_deq_bits_ops_op1),
    .io_deq_bits_ops_op2(s2_datas_io_deq_bits_ops_op2)
  );
  assign io_dmem_req_valid = io_fu_in_valid; // @[lsu.scala 100:21]
  assign io_dmem_req_bits_is_cached = io_fu_in_bits_is_cached; // @[lsu.scala 101:31]
  assign io_dmem_req_bits_addr = io_fu_in_bits_ops_op1 & 32'hfffffffc; // @[lsu.scala 102:26]
  assign io_dmem_req_bits_len = io_fu_in_bits_ops_fu_op[2:1]; // @[lsu.scala 103:26]
  assign io_dmem_req_bits_strb = _T_108[3:0]; // @[lsu.scala 106:26]
  assign io_dmem_req_bits_data = _T_95[31:0]; // @[lsu.scala 105:26]
  assign io_dmem_req_bits_func = io_fu_in_bits_ops_fu_op[3]; // @[lsu.scala 104:26]
  assign io_dmem_resp_ready = 1'h1; // @[lsu.scala 107:22]
  assign io_fu_in_ready = _T_30 | io_dmem_req_ready; // @[lsu.scala 90:18]
  assign io_fu_out_valid = io_dmem_resp_valid; // @[lsu.scala 117:19]
  assign io_fu_out_bits_v = _T_220 | _T_224; // @[lsu.scala 118:20]
  assign io_fu_out_bits_id = s2_datas_io_deq_bits_wb_id; // @[lsu.scala 120:21]
  assign io_fu_out_bits_pc = s2_datas_io_deq_bits_wb_pc; // @[lsu.scala 119:21]
  assign io_fu_out_bits_instr_op = s2_datas_io_deq_bits_wb_instr_op; // @[lsu.scala 123:24]
  assign io_fu_out_bits_instr_rs_idx = s2_datas_io_deq_bits_wb_instr_rs_idx; // @[lsu.scala 123:24]
  assign io_fu_out_bits_instr_rt_idx = s2_datas_io_deq_bits_wb_instr_rt_idx; // @[lsu.scala 123:24]
  assign io_fu_out_bits_instr_rd_idx = s2_datas_io_deq_bits_wb_instr_rd_idx; // @[lsu.scala 123:24]
  assign io_fu_out_bits_instr_shamt = s2_datas_io_deq_bits_wb_instr_shamt; // @[lsu.scala 123:24]
  assign io_fu_out_bits_instr_func = s2_datas_io_deq_bits_wb_instr_func; // @[lsu.scala 123:24]
  assign io_fu_out_bits_rd_idx = s2_datas_io_deq_bits_wb_rd_idx; // @[lsu.scala 122:25]
  assign io_fu_out_bits_wen = _T_220 | _T_224; // @[lsu.scala 121:22]
  assign io_fu_out_bits_data = _T_254[31:0]; // @[lsu.scala 128:23]
  assign io_fu_out_bits_ip7 = s2_datas_io_deq_bits_wb_ip7; // @[lsu.scala 125:22]
  assign io_fu_out_bits_is_br = s2_datas_io_deq_bits_wb_is_br; // @[lsu.scala 126:24]
  assign io_fu_out_bits_npc = s2_datas_io_deq_bits_wb_npc; // @[lsu.scala 127:22]
  assign io_working = s2_datas_io_deq_valid; // @[lsu.scala 99:14]
  assign s2_datas_clock = clock;
  assign s2_datas_reset = reset;
  assign s2_datas_io_enq_valid = io_dmem_req_ready & io_dmem_req_valid; // @[lsu.scala 96:25]
  assign s2_datas_io_enq_bits_wb_id = io_fu_in_bits_wb_id; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_pc = io_fu_in_bits_wb_pc; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_wb_npc = io_fu_in_bits_wb_npc; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_ops_fu_op = io_fu_in_bits_ops_fu_op; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_ops_op1 = io_fu_in_bits_ops_op1; // @[lsu.scala 97:24]
  assign s2_datas_io_enq_bits_ops_op2 = io_fu_in_bits_ops_op2; // @[lsu.scala 97:24]
  assign s2_datas_io_deq_ready = io_dmem_resp_ready & io_dmem_resp_valid; // @[lsu.scala 98:25]
endmodule
module MDU_Multiplier(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input  [5:0]  io_fu_in_bits_id,
  input  [4:0]  io_fu_in_bits_fu_op,
  input  [31:0] io_fu_in_bits_op1,
  input  [31:0] io_fu_in_bits_op2,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_ip7,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  output        io_fu_out_valid,
  output [5:0]  io_fu_out_bits_id,
  output [31:0] io_fu_out_bits_hi,
  output [31:0] io_fu_out_bits_lo,
  output [31:0] io_fu_out_bits_op1,
  output [4:0]  io_fu_out_bits_fu_op,
  output [7:0]  io_fu_out_bits_wb_id,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output [4:0]  io_fu_out_bits_wb_rd_idx,
  output        io_fu_out_bits_wb_ip7,
  output        io_fu_out_bits_wb_is_ds,
  output        io_fu_out_bits_wb_is_br,
  output [31:0] io_fu_out_bits_wb_npc,
  output [32:0] io_multiplier_data_a,
  output [32:0] io_multiplier_data_b,
  input  [65:0] io_multiplier_data_dout
);
  wire  _T_1 = io_fu_in_ready & io_fu_in_valid; // @[Decoupled.scala 40:37]
  reg  fu_pipePipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [5:0] fu_pipePipe_bits_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg [4:0] fu_pipePipe_bits_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg [31:0] fu_pipePipe_bits_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg [7:0] fu_pipePipe_bits_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg [31:0] fu_pipePipe_bits_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg [5:0] fu_pipePipe_bits_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg [4:0] fu_pipePipe_bits_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg [4:0] fu_pipePipe_bits_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg [4:0] fu_pipePipe_bits_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg [4:0] fu_pipePipe_bits_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg [5:0] fu_pipePipe_bits_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg [4:0] fu_pipePipe_bits_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg  fu_pipePipe_bits_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg  fu_pipePipe_bits_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg  fu_pipePipe_bits_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg [31:0] fu_pipePipe_bits_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg  fu_pipePipe_valid_1; // @[Valid.scala 117:22]
  reg [31:0] _RAND_17;
  reg [5:0] fu_pipePipe_bits_1_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg [4:0] fu_pipePipe_bits_1_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg [31:0] fu_pipePipe_bits_1_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg [7:0] fu_pipePipe_bits_1_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg [31:0] fu_pipePipe_bits_1_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg [5:0] fu_pipePipe_bits_1_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg [4:0] fu_pipePipe_bits_1_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg [4:0] fu_pipePipe_bits_1_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg [4:0] fu_pipePipe_bits_1_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg [4:0] fu_pipePipe_bits_1_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg [5:0] fu_pipePipe_bits_1_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg [4:0] fu_pipePipe_bits_1_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  fu_pipePipe_bits_1_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg  fu_pipePipe_bits_1_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg  fu_pipePipe_bits_1_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg [31:0] fu_pipePipe_bits_1_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg  fu_pipePipe_valid_2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_34;
  reg [5:0] fu_pipePipe_bits_2_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg [4:0] fu_pipePipe_bits_2_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg [31:0] fu_pipePipe_bits_2_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg [7:0] fu_pipePipe_bits_2_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg [31:0] fu_pipePipe_bits_2_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg [5:0] fu_pipePipe_bits_2_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg [4:0] fu_pipePipe_bits_2_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg [4:0] fu_pipePipe_bits_2_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg [4:0] fu_pipePipe_bits_2_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg [4:0] fu_pipePipe_bits_2_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg [5:0] fu_pipePipe_bits_2_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg [4:0] fu_pipePipe_bits_2_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg  fu_pipePipe_bits_2_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg  fu_pipePipe_bits_2_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg  fu_pipePipe_bits_2_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg [31:0] fu_pipePipe_bits_2_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg  fu_pipePipe_valid_3; // @[Valid.scala 117:22]
  reg [31:0] _RAND_51;
  reg [5:0] fu_pipePipe_bits_3_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg [4:0] fu_pipePipe_bits_3_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg [31:0] fu_pipePipe_bits_3_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg [7:0] fu_pipePipe_bits_3_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg [31:0] fu_pipePipe_bits_3_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg [5:0] fu_pipePipe_bits_3_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg [4:0] fu_pipePipe_bits_3_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg [4:0] fu_pipePipe_bits_3_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg [4:0] fu_pipePipe_bits_3_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg [4:0] fu_pipePipe_bits_3_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg [5:0] fu_pipePipe_bits_3_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg [4:0] fu_pipePipe_bits_3_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg  fu_pipePipe_bits_3_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg  fu_pipePipe_bits_3_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg  fu_pipePipe_bits_3_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg [31:0] fu_pipePipe_bits_3_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg  fu_pipePipe_valid_4; // @[Valid.scala 117:22]
  reg [31:0] _RAND_68;
  reg [5:0] fu_pipePipe_bits_4_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg [4:0] fu_pipePipe_bits_4_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg [31:0] fu_pipePipe_bits_4_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg [7:0] fu_pipePipe_bits_4_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg [31:0] fu_pipePipe_bits_4_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg [5:0] fu_pipePipe_bits_4_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg [4:0] fu_pipePipe_bits_4_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg [4:0] fu_pipePipe_bits_4_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg [4:0] fu_pipePipe_bits_4_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg [4:0] fu_pipePipe_bits_4_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg [5:0] fu_pipePipe_bits_4_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg [4:0] fu_pipePipe_bits_4_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg  fu_pipePipe_bits_4_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg  fu_pipePipe_bits_4_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg  fu_pipePipe_bits_4_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg [31:0] fu_pipePipe_bits_4_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg  fu_pipePipe_valid_5; // @[Valid.scala 117:22]
  reg [31:0] _RAND_85;
  reg [5:0] fu_pipePipe_bits_5_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg [4:0] fu_pipePipe_bits_5_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg [31:0] fu_pipePipe_bits_5_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg [7:0] fu_pipePipe_bits_5_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg [31:0] fu_pipePipe_bits_5_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg [5:0] fu_pipePipe_bits_5_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg [4:0] fu_pipePipe_bits_5_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg [4:0] fu_pipePipe_bits_5_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg [4:0] fu_pipePipe_bits_5_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg [4:0] fu_pipePipe_bits_5_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg [5:0] fu_pipePipe_bits_5_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg [4:0] fu_pipePipe_bits_5_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg  fu_pipePipe_bits_5_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg  fu_pipePipe_bits_5_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg  fu_pipePipe_bits_5_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg [31:0] fu_pipePipe_bits_5_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg  fu_pipePipe_valid_6; // @[Valid.scala 117:22]
  reg [31:0] _RAND_102;
  reg [5:0] fu_pipePipe_bits_6_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg [4:0] fu_pipePipe_bits_6_fu_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg [31:0] fu_pipePipe_bits_6_op1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg [7:0] fu_pipePipe_bits_6_wb_id; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg [31:0] fu_pipePipe_bits_6_wb_pc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg [5:0] fu_pipePipe_bits_6_wb_instr_op; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg [4:0] fu_pipePipe_bits_6_wb_instr_rs_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg [4:0] fu_pipePipe_bits_6_wb_instr_rt_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg [4:0] fu_pipePipe_bits_6_wb_instr_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg [4:0] fu_pipePipe_bits_6_wb_instr_shamt; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg [5:0] fu_pipePipe_bits_6_wb_instr_func; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg [4:0] fu_pipePipe_bits_6_wb_rd_idx; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg  fu_pipePipe_bits_6_wb_ip7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg  fu_pipePipe_bits_6_wb_is_ds; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg  fu_pipePipe_bits_6_wb_is_br; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg [31:0] fu_pipePipe_bits_6_wb_npc; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  wire  _T_2 = io_fu_in_bits_fu_op == 5'hb; // @[mdu.scala 57:45]
  wire [31:0] _T_4 = io_fu_in_bits_op1; // @[mdu.scala 58:17]
  wire [32:0] _T_5 = {{1{_T_4[31]}},_T_4}; // @[mdu.scala 58:30]
  wire [32:0] _T_6 = {{1'd0}, io_fu_in_bits_op1}; // @[mdu.scala 59:17 mdu.scala 59:17]
  wire [31:0] _T_10 = io_fu_in_bits_op2; // @[mdu.scala 61:17]
  wire [32:0] _T_11 = {{1{_T_10[31]}},_T_10}; // @[mdu.scala 61:30]
  wire [32:0] _T_12 = {{1'd0}, io_fu_in_bits_op2}; // @[mdu.scala 62:17 mdu.scala 62:17]
  assign io_fu_in_ready = 1'h1; // @[mdu.scala 64:18]
  assign io_fu_out_valid = fu_pipePipe_valid_6; // @[mdu.scala 65:19]
  assign io_fu_out_bits_id = fu_pipePipe_bits_6_id; // @[mdu.scala 68:21]
  assign io_fu_out_bits_hi = io_multiplier_data_dout[63:32]; // @[mdu.scala 70:21]
  assign io_fu_out_bits_lo = io_multiplier_data_dout[31:0]; // @[mdu.scala 71:21]
  assign io_fu_out_bits_op1 = fu_pipePipe_bits_6_op1; // @[mdu.scala 69:22]
  assign io_fu_out_bits_fu_op = fu_pipePipe_bits_6_fu_op; // @[mdu.scala 66:24]
  assign io_fu_out_bits_wb_id = fu_pipePipe_bits_6_wb_id; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_pc = fu_pipePipe_bits_6_wb_pc; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_instr_op = fu_pipePipe_bits_6_wb_instr_op; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_instr_rs_idx = fu_pipePipe_bits_6_wb_instr_rs_idx; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_instr_rt_idx = fu_pipePipe_bits_6_wb_instr_rt_idx; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_instr_rd_idx = fu_pipePipe_bits_6_wb_instr_rd_idx; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_instr_shamt = fu_pipePipe_bits_6_wb_instr_shamt; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_instr_func = fu_pipePipe_bits_6_wb_instr_func; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_rd_idx = fu_pipePipe_bits_6_wb_rd_idx; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_ip7 = fu_pipePipe_bits_6_wb_ip7; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_is_ds = fu_pipePipe_bits_6_wb_is_ds; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_is_br = fu_pipePipe_bits_6_wb_is_br; // @[mdu.scala 67:21]
  assign io_fu_out_bits_wb_npc = fu_pipePipe_bits_6_wb_npc; // @[mdu.scala 67:21]
  assign io_multiplier_data_a = _T_2 ? _T_5 : _T_6; // @[mdu.scala 57:24]
  assign io_multiplier_data_b = _T_2 ? _T_11 : _T_12; // @[mdu.scala 60:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fu_pipePipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fu_pipePipe_bits_id = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  fu_pipePipe_bits_fu_op = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fu_pipePipe_bits_op1 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_id = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_instr_op = _RAND_6[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_instr_rs_idx = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_instr_rt_idx = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_instr_rd_idx = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_instr_shamt = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_instr_func = _RAND_11[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_rd_idx = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_ip7 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_is_ds = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_is_br = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  fu_pipePipe_bits_wb_npc = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  fu_pipePipe_valid_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  fu_pipePipe_bits_1_id = _RAND_18[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  fu_pipePipe_bits_1_fu_op = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  fu_pipePipe_bits_1_op1 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_id = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_pc = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_instr_op = _RAND_23[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_instr_rs_idx = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_instr_rt_idx = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_instr_rd_idx = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_instr_shamt = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_instr_func = _RAND_28[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_rd_idx = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_ip7 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_is_ds = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_is_br = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  fu_pipePipe_bits_1_wb_npc = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  fu_pipePipe_valid_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  fu_pipePipe_bits_2_id = _RAND_35[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  fu_pipePipe_bits_2_fu_op = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  fu_pipePipe_bits_2_op1 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_id = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_pc = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_instr_op = _RAND_40[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_instr_rs_idx = _RAND_41[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_instr_rt_idx = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_instr_rd_idx = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_instr_shamt = _RAND_44[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_instr_func = _RAND_45[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_rd_idx = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_ip7 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_is_ds = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_is_br = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  fu_pipePipe_bits_2_wb_npc = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  fu_pipePipe_valid_3 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  fu_pipePipe_bits_3_id = _RAND_52[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  fu_pipePipe_bits_3_fu_op = _RAND_53[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  fu_pipePipe_bits_3_op1 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_id = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_pc = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_instr_op = _RAND_57[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_instr_rs_idx = _RAND_58[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_instr_rt_idx = _RAND_59[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_instr_rd_idx = _RAND_60[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_instr_shamt = _RAND_61[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_instr_func = _RAND_62[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_rd_idx = _RAND_63[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_ip7 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_is_ds = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_is_br = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  fu_pipePipe_bits_3_wb_npc = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  fu_pipePipe_valid_4 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  fu_pipePipe_bits_4_id = _RAND_69[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  fu_pipePipe_bits_4_fu_op = _RAND_70[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  fu_pipePipe_bits_4_op1 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_id = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_pc = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_instr_op = _RAND_74[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_instr_rs_idx = _RAND_75[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_instr_rt_idx = _RAND_76[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_instr_rd_idx = _RAND_77[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_instr_shamt = _RAND_78[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_instr_func = _RAND_79[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_rd_idx = _RAND_80[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_ip7 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_is_ds = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_is_br = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  fu_pipePipe_bits_4_wb_npc = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  fu_pipePipe_valid_5 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  fu_pipePipe_bits_5_id = _RAND_86[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  fu_pipePipe_bits_5_fu_op = _RAND_87[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  fu_pipePipe_bits_5_op1 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_id = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_pc = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_instr_op = _RAND_91[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_instr_rs_idx = _RAND_92[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_instr_rt_idx = _RAND_93[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_instr_rd_idx = _RAND_94[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_instr_shamt = _RAND_95[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_instr_func = _RAND_96[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_rd_idx = _RAND_97[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_ip7 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_is_ds = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_is_br = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  fu_pipePipe_bits_5_wb_npc = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  fu_pipePipe_valid_6 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  fu_pipePipe_bits_6_id = _RAND_103[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  fu_pipePipe_bits_6_fu_op = _RAND_104[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  fu_pipePipe_bits_6_op1 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_id = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_pc = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_instr_op = _RAND_108[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_instr_rs_idx = _RAND_109[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_instr_rt_idx = _RAND_110[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_instr_rd_idx = _RAND_111[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_instr_shamt = _RAND_112[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_instr_func = _RAND_113[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_rd_idx = _RAND_114[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_ip7 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_is_ds = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_is_br = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  fu_pipePipe_bits_6_wb_npc = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fu_pipePipe_valid <= 1'h0;
    end else begin
      fu_pipePipe_valid <= _T_1;
    end
    if (_T_1) begin
      fu_pipePipe_bits_id <= io_fu_in_bits_id;
    end
    if (_T_1) begin
      fu_pipePipe_bits_fu_op <= io_fu_in_bits_fu_op;
    end
    if (_T_1) begin
      fu_pipePipe_bits_op1 <= io_fu_in_bits_op1;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_id <= io_fu_in_bits_wb_id;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_pc <= io_fu_in_bits_wb_pc;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_instr_op <= io_fu_in_bits_wb_instr_op;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_instr_rs_idx <= io_fu_in_bits_wb_instr_rs_idx;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_instr_rt_idx <= io_fu_in_bits_wb_instr_rt_idx;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_instr_rd_idx <= io_fu_in_bits_wb_instr_rd_idx;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_instr_shamt <= io_fu_in_bits_wb_instr_shamt;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_instr_func <= io_fu_in_bits_wb_instr_func;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_rd_idx <= io_fu_in_bits_wb_rd_idx;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_ip7 <= io_fu_in_bits_wb_ip7;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_is_ds <= io_fu_in_bits_wb_is_ds;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_is_br <= io_fu_in_bits_wb_is_br;
    end
    if (_T_1) begin
      fu_pipePipe_bits_wb_npc <= io_fu_in_bits_wb_npc;
    end
    if (reset) begin
      fu_pipePipe_valid_1 <= 1'h0;
    end else begin
      fu_pipePipe_valid_1 <= fu_pipePipe_valid;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_id <= fu_pipePipe_bits_id;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_fu_op <= fu_pipePipe_bits_fu_op;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_op1 <= fu_pipePipe_bits_op1;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_id <= fu_pipePipe_bits_wb_id;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_pc <= fu_pipePipe_bits_wb_pc;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_instr_op <= fu_pipePipe_bits_wb_instr_op;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_instr_rs_idx <= fu_pipePipe_bits_wb_instr_rs_idx;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_instr_rt_idx <= fu_pipePipe_bits_wb_instr_rt_idx;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_instr_rd_idx <= fu_pipePipe_bits_wb_instr_rd_idx;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_instr_shamt <= fu_pipePipe_bits_wb_instr_shamt;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_instr_func <= fu_pipePipe_bits_wb_instr_func;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_rd_idx <= fu_pipePipe_bits_wb_rd_idx;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_ip7 <= fu_pipePipe_bits_wb_ip7;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_is_ds <= fu_pipePipe_bits_wb_is_ds;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_is_br <= fu_pipePipe_bits_wb_is_br;
    end
    if (fu_pipePipe_valid) begin
      fu_pipePipe_bits_1_wb_npc <= fu_pipePipe_bits_wb_npc;
    end
    if (reset) begin
      fu_pipePipe_valid_2 <= 1'h0;
    end else begin
      fu_pipePipe_valid_2 <= fu_pipePipe_valid_1;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_id <= fu_pipePipe_bits_1_id;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_fu_op <= fu_pipePipe_bits_1_fu_op;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_op1 <= fu_pipePipe_bits_1_op1;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_id <= fu_pipePipe_bits_1_wb_id;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_pc <= fu_pipePipe_bits_1_wb_pc;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_instr_op <= fu_pipePipe_bits_1_wb_instr_op;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_instr_rs_idx <= fu_pipePipe_bits_1_wb_instr_rs_idx;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_instr_rt_idx <= fu_pipePipe_bits_1_wb_instr_rt_idx;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_instr_rd_idx <= fu_pipePipe_bits_1_wb_instr_rd_idx;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_instr_shamt <= fu_pipePipe_bits_1_wb_instr_shamt;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_instr_func <= fu_pipePipe_bits_1_wb_instr_func;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_rd_idx <= fu_pipePipe_bits_1_wb_rd_idx;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_ip7 <= fu_pipePipe_bits_1_wb_ip7;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_is_ds <= fu_pipePipe_bits_1_wb_is_ds;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_is_br <= fu_pipePipe_bits_1_wb_is_br;
    end
    if (fu_pipePipe_valid_1) begin
      fu_pipePipe_bits_2_wb_npc <= fu_pipePipe_bits_1_wb_npc;
    end
    if (reset) begin
      fu_pipePipe_valid_3 <= 1'h0;
    end else begin
      fu_pipePipe_valid_3 <= fu_pipePipe_valid_2;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_id <= fu_pipePipe_bits_2_id;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_fu_op <= fu_pipePipe_bits_2_fu_op;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_op1 <= fu_pipePipe_bits_2_op1;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_id <= fu_pipePipe_bits_2_wb_id;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_pc <= fu_pipePipe_bits_2_wb_pc;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_instr_op <= fu_pipePipe_bits_2_wb_instr_op;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_instr_rs_idx <= fu_pipePipe_bits_2_wb_instr_rs_idx;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_instr_rt_idx <= fu_pipePipe_bits_2_wb_instr_rt_idx;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_instr_rd_idx <= fu_pipePipe_bits_2_wb_instr_rd_idx;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_instr_shamt <= fu_pipePipe_bits_2_wb_instr_shamt;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_instr_func <= fu_pipePipe_bits_2_wb_instr_func;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_rd_idx <= fu_pipePipe_bits_2_wb_rd_idx;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_ip7 <= fu_pipePipe_bits_2_wb_ip7;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_is_ds <= fu_pipePipe_bits_2_wb_is_ds;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_is_br <= fu_pipePipe_bits_2_wb_is_br;
    end
    if (fu_pipePipe_valid_2) begin
      fu_pipePipe_bits_3_wb_npc <= fu_pipePipe_bits_2_wb_npc;
    end
    if (reset) begin
      fu_pipePipe_valid_4 <= 1'h0;
    end else begin
      fu_pipePipe_valid_4 <= fu_pipePipe_valid_3;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_id <= fu_pipePipe_bits_3_id;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_fu_op <= fu_pipePipe_bits_3_fu_op;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_op1 <= fu_pipePipe_bits_3_op1;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_id <= fu_pipePipe_bits_3_wb_id;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_pc <= fu_pipePipe_bits_3_wb_pc;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_instr_op <= fu_pipePipe_bits_3_wb_instr_op;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_instr_rs_idx <= fu_pipePipe_bits_3_wb_instr_rs_idx;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_instr_rt_idx <= fu_pipePipe_bits_3_wb_instr_rt_idx;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_instr_rd_idx <= fu_pipePipe_bits_3_wb_instr_rd_idx;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_instr_shamt <= fu_pipePipe_bits_3_wb_instr_shamt;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_instr_func <= fu_pipePipe_bits_3_wb_instr_func;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_rd_idx <= fu_pipePipe_bits_3_wb_rd_idx;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_ip7 <= fu_pipePipe_bits_3_wb_ip7;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_is_ds <= fu_pipePipe_bits_3_wb_is_ds;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_is_br <= fu_pipePipe_bits_3_wb_is_br;
    end
    if (fu_pipePipe_valid_3) begin
      fu_pipePipe_bits_4_wb_npc <= fu_pipePipe_bits_3_wb_npc;
    end
    if (reset) begin
      fu_pipePipe_valid_5 <= 1'h0;
    end else begin
      fu_pipePipe_valid_5 <= fu_pipePipe_valid_4;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_id <= fu_pipePipe_bits_4_id;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_fu_op <= fu_pipePipe_bits_4_fu_op;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_op1 <= fu_pipePipe_bits_4_op1;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_id <= fu_pipePipe_bits_4_wb_id;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_pc <= fu_pipePipe_bits_4_wb_pc;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_instr_op <= fu_pipePipe_bits_4_wb_instr_op;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_instr_rs_idx <= fu_pipePipe_bits_4_wb_instr_rs_idx;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_instr_rt_idx <= fu_pipePipe_bits_4_wb_instr_rt_idx;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_instr_rd_idx <= fu_pipePipe_bits_4_wb_instr_rd_idx;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_instr_shamt <= fu_pipePipe_bits_4_wb_instr_shamt;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_instr_func <= fu_pipePipe_bits_4_wb_instr_func;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_rd_idx <= fu_pipePipe_bits_4_wb_rd_idx;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_ip7 <= fu_pipePipe_bits_4_wb_ip7;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_is_ds <= fu_pipePipe_bits_4_wb_is_ds;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_is_br <= fu_pipePipe_bits_4_wb_is_br;
    end
    if (fu_pipePipe_valid_4) begin
      fu_pipePipe_bits_5_wb_npc <= fu_pipePipe_bits_4_wb_npc;
    end
    if (reset) begin
      fu_pipePipe_valid_6 <= 1'h0;
    end else begin
      fu_pipePipe_valid_6 <= fu_pipePipe_valid_5;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_id <= fu_pipePipe_bits_5_id;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_fu_op <= fu_pipePipe_bits_5_fu_op;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_op1 <= fu_pipePipe_bits_5_op1;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_id <= fu_pipePipe_bits_5_wb_id;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_pc <= fu_pipePipe_bits_5_wb_pc;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_instr_op <= fu_pipePipe_bits_5_wb_instr_op;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_instr_rs_idx <= fu_pipePipe_bits_5_wb_instr_rs_idx;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_instr_rt_idx <= fu_pipePipe_bits_5_wb_instr_rt_idx;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_instr_rd_idx <= fu_pipePipe_bits_5_wb_instr_rd_idx;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_instr_shamt <= fu_pipePipe_bits_5_wb_instr_shamt;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_instr_func <= fu_pipePipe_bits_5_wb_instr_func;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_rd_idx <= fu_pipePipe_bits_5_wb_rd_idx;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_ip7 <= fu_pipePipe_bits_5_wb_ip7;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_is_ds <= fu_pipePipe_bits_5_wb_is_ds;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_is_br <= fu_pipePipe_bits_5_wb_is_br;
    end
    if (fu_pipePipe_valid_5) begin
      fu_pipePipe_bits_6_wb_npc <= fu_pipePipe_bits_5_wb_npc;
    end
  end
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [5:0]  io_enq_bits_id,
  input  [4:0]  io_enq_bits_fu_op,
  input  [31:0] io_enq_bits_op1,
  input  [7:0]  io_enq_bits_wb_id,
  input  [31:0] io_enq_bits_wb_pc,
  input  [5:0]  io_enq_bits_wb_instr_op,
  input  [4:0]  io_enq_bits_wb_instr_rs_idx,
  input  [4:0]  io_enq_bits_wb_instr_rt_idx,
  input  [4:0]  io_enq_bits_wb_instr_rd_idx,
  input  [4:0]  io_enq_bits_wb_instr_shamt,
  input  [5:0]  io_enq_bits_wb_instr_func,
  input  [4:0]  io_enq_bits_wb_rd_idx,
  input         io_enq_bits_wb_ip7,
  input         io_enq_bits_wb_is_ds,
  input         io_enq_bits_wb_is_br,
  input  [31:0] io_enq_bits_wb_npc,
  input         io_deq_ready,
  output        io_deq_valid,
  output [5:0]  io_deq_bits_id,
  output [4:0]  io_deq_bits_fu_op,
  output [31:0] io_deq_bits_op1,
  output [7:0]  io_deq_bits_wb_id,
  output [31:0] io_deq_bits_wb_pc,
  output [5:0]  io_deq_bits_wb_instr_op,
  output [4:0]  io_deq_bits_wb_instr_rs_idx,
  output [4:0]  io_deq_bits_wb_instr_rt_idx,
  output [4:0]  io_deq_bits_wb_instr_rd_idx,
  output [4:0]  io_deq_bits_wb_instr_shamt,
  output [5:0]  io_deq_bits_wb_instr_func,
  output [4:0]  io_deq_bits_wb_rd_idx,
  output        io_deq_bits_wb_ip7,
  output        io_deq_bits_wb_is_ds,
  output        io_deq_bits_wb_is_br,
  output [31:0] io_deq_bits_wb_npc
);
  reg [5:0] _T_id [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_0;
  wire [5:0] _T_id__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_id__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_1;
  wire [5:0] _T_id__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_id__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_id__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_fu_op [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_2;
  wire [4:0] _T_fu_op__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_fu_op__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_3;
  wire [4:0] _T_fu_op__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_fu_op__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_fu_op__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_fu_op__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_op1 [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_4;
  wire [31:0] _T_op1__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_op1__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_5;
  wire [31:0] _T_op1__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_op1__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_op1__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_op1__T_10_en; // @[Decoupled.scala 218:24]
  reg [7:0] _T_wb_id [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_6;
  wire [7:0] _T_wb_id__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_id__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_7;
  wire [7:0] _T_wb_id__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_id__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_id__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_id__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_wb_pc [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_8;
  wire [31:0] _T_wb_pc__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_pc__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_9;
  wire [31:0] _T_wb_pc__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_pc__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_pc__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_pc__T_10_en; // @[Decoupled.scala 218:24]
  reg [5:0] _T_wb_instr_op [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_10;
  wire [5:0] _T_wb_instr_op__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_op__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_11;
  wire [5:0] _T_wb_instr_op__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_op__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_op__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_op__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_rs_idx [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_12;
  wire [4:0] _T_wb_instr_rs_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_rs_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_13;
  wire [4:0] _T_wb_instr_rs_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_rs_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rs_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rs_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_rt_idx [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_14;
  wire [4:0] _T_wb_instr_rt_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_rt_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_15;
  wire [4:0] _T_wb_instr_rt_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_rt_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rt_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rt_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_rd_idx [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_16;
  wire [4:0] _T_wb_instr_rd_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_rd_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_17;
  wire [4:0] _T_wb_instr_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_rd_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rd_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_rd_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_instr_shamt [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_18;
  wire [4:0] _T_wb_instr_shamt__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_shamt__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_19;
  wire [4:0] _T_wb_instr_shamt__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_shamt__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_shamt__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_shamt__T_10_en; // @[Decoupled.scala 218:24]
  reg [5:0] _T_wb_instr_func [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_20;
  wire [5:0] _T_wb_instr_func__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_func__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_21;
  wire [5:0] _T_wb_instr_func__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_instr_func__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_func__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_instr_func__T_10_en; // @[Decoupled.scala 218:24]
  reg [4:0] _T_wb_rd_idx [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_22;
  wire [4:0] _T_wb_rd_idx__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_rd_idx__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_23;
  wire [4:0] _T_wb_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_rd_idx__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_rd_idx__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_rd_idx__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_wb_ip7 [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_24;
  wire  _T_wb_ip7__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_ip7__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_25;
  wire  _T_wb_ip7__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_ip7__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_ip7__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_ip7__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_wb_is_ds [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_26;
  wire  _T_wb_is_ds__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_is_ds__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_27;
  wire  _T_wb_is_ds__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_is_ds__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_is_ds__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_is_ds__T_10_en; // @[Decoupled.scala 218:24]
  reg  _T_wb_is_br [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_28;
  wire  _T_wb_is_br__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_is_br__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_29;
  wire  _T_wb_is_br__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_is_br__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_is_br__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_is_br__T_10_en; // @[Decoupled.scala 218:24]
  reg [31:0] _T_wb_npc [0:44]; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_30;
  wire [31:0] _T_wb_npc__T_18_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_npc__T_18_addr; // @[Decoupled.scala 218:24]
  reg [31:0] _RAND_31;
  wire [31:0] _T_wb_npc__T_10_data; // @[Decoupled.scala 218:24]
  wire [5:0] _T_wb_npc__T_10_addr; // @[Decoupled.scala 218:24]
  wire  _T_wb_npc__T_10_mask; // @[Decoupled.scala 218:24]
  wire  _T_wb_npc__T_10_en; // @[Decoupled.scala 218:24]
  reg [5:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_32;
  reg [5:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_33;
  reg  _T_1; // @[Decoupled.scala 221:35]
  reg [31:0] _RAND_34;
  wire  _T_2 = value == value_1; // @[Decoupled.scala 223:41]
  wire  _T_3 = ~_T_1; // @[Decoupled.scala 224:36]
  wire  _T_4 = _T_2 & _T_3; // @[Decoupled.scala 224:33]
  wire  _T_5 = _T_2 & _T_1; // @[Decoupled.scala 225:32]
  wire  _T_6 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_8 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = value == 6'h2c; // @[Counter.scala 38:24]
  wire [5:0] _T_12 = value + 6'h1; // @[Counter.scala 39:22]
  wire  wrap_1 = value_1 == 6'h2c; // @[Counter.scala 38:24]
  wire [5:0] _T_14 = value_1 + 6'h1; // @[Counter.scala 39:22]
  wire  _T_15 = _T_6 != _T_8; // @[Decoupled.scala 236:16]
  assign _T_id__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_id__T_18_data = _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_id__T_18_data = _T_id__T_18_addr >= 6'h2d ? _RAND_1[5:0] : _T_id[_T_id__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_id__T_10_data = io_enq_bits_id;
  assign _T_id__T_10_addr = value;
  assign _T_id__T_10_mask = 1'h1;
  assign _T_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_fu_op__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_fu_op__T_18_data = _T_fu_op[_T_fu_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_fu_op__T_18_data = _T_fu_op__T_18_addr >= 6'h2d ? _RAND_3[4:0] : _T_fu_op[_T_fu_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_fu_op__T_10_data = io_enq_bits_fu_op;
  assign _T_fu_op__T_10_addr = value;
  assign _T_fu_op__T_10_mask = 1'h1;
  assign _T_fu_op__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_op1__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_op1__T_18_data = _T_op1[_T_op1__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_op1__T_18_data = _T_op1__T_18_addr >= 6'h2d ? _RAND_5[31:0] : _T_op1[_T_op1__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_op1__T_10_data = io_enq_bits_op1;
  assign _T_op1__T_10_addr = value;
  assign _T_op1__T_10_mask = 1'h1;
  assign _T_op1__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_id__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_id__T_18_data = _T_wb_id[_T_wb_id__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_id__T_18_data = _T_wb_id__T_18_addr >= 6'h2d ? _RAND_7[7:0] : _T_wb_id[_T_wb_id__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_id__T_10_data = io_enq_bits_wb_id;
  assign _T_wb_id__T_10_addr = value;
  assign _T_wb_id__T_10_mask = 1'h1;
  assign _T_wb_id__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_pc__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_pc__T_18_data = _T_wb_pc[_T_wb_pc__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_pc__T_18_data = _T_wb_pc__T_18_addr >= 6'h2d ? _RAND_9[31:0] : _T_wb_pc[_T_wb_pc__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_pc__T_10_data = io_enq_bits_wb_pc;
  assign _T_wb_pc__T_10_addr = value;
  assign _T_wb_pc__T_10_mask = 1'h1;
  assign _T_wb_pc__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_op__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_op__T_18_data = _T_wb_instr_op[_T_wb_instr_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_op__T_18_data = _T_wb_instr_op__T_18_addr >= 6'h2d ? _RAND_11[5:0] : _T_wb_instr_op[_T_wb_instr_op__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_op__T_10_data = io_enq_bits_wb_instr_op;
  assign _T_wb_instr_op__T_10_addr = value;
  assign _T_wb_instr_op__T_10_mask = 1'h1;
  assign _T_wb_instr_op__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_rs_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rs_idx__T_18_data = _T_wb_instr_rs_idx[_T_wb_instr_rs_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_rs_idx__T_18_data = _T_wb_instr_rs_idx__T_18_addr >= 6'h2d ? _RAND_13[4:0] : _T_wb_instr_rs_idx[_T_wb_instr_rs_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rs_idx__T_10_data = io_enq_bits_wb_instr_rs_idx;
  assign _T_wb_instr_rs_idx__T_10_addr = value;
  assign _T_wb_instr_rs_idx__T_10_mask = 1'h1;
  assign _T_wb_instr_rs_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_rt_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rt_idx__T_18_data = _T_wb_instr_rt_idx[_T_wb_instr_rt_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_rt_idx__T_18_data = _T_wb_instr_rt_idx__T_18_addr >= 6'h2d ? _RAND_15[4:0] : _T_wb_instr_rt_idx[_T_wb_instr_rt_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rt_idx__T_10_data = io_enq_bits_wb_instr_rt_idx;
  assign _T_wb_instr_rt_idx__T_10_addr = value;
  assign _T_wb_instr_rt_idx__T_10_mask = 1'h1;
  assign _T_wb_instr_rt_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_rd_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rd_idx__T_18_data = _T_wb_instr_rd_idx[_T_wb_instr_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_rd_idx__T_18_data = _T_wb_instr_rd_idx__T_18_addr >= 6'h2d ? _RAND_17[4:0] : _T_wb_instr_rd_idx[_T_wb_instr_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_rd_idx__T_10_data = io_enq_bits_wb_instr_rd_idx;
  assign _T_wb_instr_rd_idx__T_10_addr = value;
  assign _T_wb_instr_rd_idx__T_10_mask = 1'h1;
  assign _T_wb_instr_rd_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_shamt__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_shamt__T_18_data = _T_wb_instr_shamt[_T_wb_instr_shamt__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_shamt__T_18_data = _T_wb_instr_shamt__T_18_addr >= 6'h2d ? _RAND_19[4:0] : _T_wb_instr_shamt[_T_wb_instr_shamt__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_shamt__T_10_data = io_enq_bits_wb_instr_shamt;
  assign _T_wb_instr_shamt__T_10_addr = value;
  assign _T_wb_instr_shamt__T_10_mask = 1'h1;
  assign _T_wb_instr_shamt__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_instr_func__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_func__T_18_data = _T_wb_instr_func[_T_wb_instr_func__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_instr_func__T_18_data = _T_wb_instr_func__T_18_addr >= 6'h2d ? _RAND_21[5:0] : _T_wb_instr_func[_T_wb_instr_func__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_instr_func__T_10_data = io_enq_bits_wb_instr_func;
  assign _T_wb_instr_func__T_10_addr = value;
  assign _T_wb_instr_func__T_10_mask = 1'h1;
  assign _T_wb_instr_func__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_rd_idx__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_rd_idx__T_18_data = _T_wb_rd_idx[_T_wb_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_rd_idx__T_18_data = _T_wb_rd_idx__T_18_addr >= 6'h2d ? _RAND_23[4:0] : _T_wb_rd_idx[_T_wb_rd_idx__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_rd_idx__T_10_data = io_enq_bits_wb_rd_idx;
  assign _T_wb_rd_idx__T_10_addr = value;
  assign _T_wb_rd_idx__T_10_mask = 1'h1;
  assign _T_wb_rd_idx__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_ip7__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_ip7__T_18_data = _T_wb_ip7[_T_wb_ip7__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_ip7__T_18_data = _T_wb_ip7__T_18_addr >= 6'h2d ? _RAND_25[0:0] : _T_wb_ip7[_T_wb_ip7__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_ip7__T_10_data = io_enq_bits_wb_ip7;
  assign _T_wb_ip7__T_10_addr = value;
  assign _T_wb_ip7__T_10_mask = 1'h1;
  assign _T_wb_ip7__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_is_ds__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_is_ds__T_18_data = _T_wb_is_ds[_T_wb_is_ds__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_is_ds__T_18_data = _T_wb_is_ds__T_18_addr >= 6'h2d ? _RAND_27[0:0] : _T_wb_is_ds[_T_wb_is_ds__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_is_ds__T_10_data = io_enq_bits_wb_is_ds;
  assign _T_wb_is_ds__T_10_addr = value;
  assign _T_wb_is_ds__T_10_mask = 1'h1;
  assign _T_wb_is_ds__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_is_br__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_is_br__T_18_data = _T_wb_is_br[_T_wb_is_br__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_is_br__T_18_data = _T_wb_is_br__T_18_addr >= 6'h2d ? _RAND_29[0:0] : _T_wb_is_br[_T_wb_is_br__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_is_br__T_10_data = io_enq_bits_wb_is_br;
  assign _T_wb_is_br__T_10_addr = value;
  assign _T_wb_is_br__T_10_mask = 1'h1;
  assign _T_wb_is_br__T_10_en = io_enq_ready & io_enq_valid;
  assign _T_wb_npc__T_18_addr = value_1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_npc__T_18_data = _T_wb_npc[_T_wb_npc__T_18_addr]; // @[Decoupled.scala 218:24]
  `else
  assign _T_wb_npc__T_18_data = _T_wb_npc__T_18_addr >= 6'h2d ? _RAND_31[31:0] : _T_wb_npc[_T_wb_npc__T_18_addr]; // @[Decoupled.scala 218:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_wb_npc__T_10_data = io_enq_bits_wb_npc;
  assign _T_wb_npc__T_10_addr = value;
  assign _T_wb_npc__T_10_mask = 1'h1;
  assign _T_wb_npc__T_10_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_5; // @[Decoupled.scala 241:16]
  assign io_deq_valid = ~_T_4; // @[Decoupled.scala 240:16]
  assign io_deq_bits_id = _T_id__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_fu_op = _T_fu_op__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_op1 = _T_op1__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_id = _T_wb_id__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_pc = _T_wb_pc__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_op = _T_wb_instr_op__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_rs_idx = _T_wb_instr_rs_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_rt_idx = _T_wb_instr_rt_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_rd_idx = _T_wb_instr_rd_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_shamt = _T_wb_instr_shamt__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_instr_func = _T_wb_instr_func__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_rd_idx = _T_wb_rd_idx__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_ip7 = _T_wb_ip7__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_is_ds = _T_wb_is_ds__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_is_br = _T_wb_is_br__T_18_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_wb_npc = _T_wb_npc__T_18_data; // @[Decoupled.scala 242:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_id[initvar] = _RAND_0[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_fu_op[initvar] = _RAND_2[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_op1[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_id[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_pc[initvar] = _RAND_8[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_instr_op[initvar] = _RAND_10[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_instr_rs_idx[initvar] = _RAND_12[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_instr_rt_idx[initvar] = _RAND_14[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_instr_rd_idx[initvar] = _RAND_16[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  _RAND_18 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_instr_shamt[initvar] = _RAND_18[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_19 = {1{`RANDOM}};
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_instr_func[initvar] = _RAND_20[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  _RAND_22 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_rd_idx[initvar] = _RAND_22[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_23 = {1{`RANDOM}};
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_ip7[initvar] = _RAND_24[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  _RAND_26 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_is_ds[initvar] = _RAND_26[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_27 = {1{`RANDOM}};
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_is_br[initvar] = _RAND_28[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  _RAND_30 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 45; initvar = initvar+1)
    _T_wb_npc[initvar] = _RAND_30[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_31 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  value = _RAND_32[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  value_1 = _RAND_33[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_1 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_id__T_10_en & _T_id__T_10_mask) begin
      _T_id[_T_id__T_10_addr] <= _T_id__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_fu_op__T_10_en & _T_fu_op__T_10_mask) begin
      _T_fu_op[_T_fu_op__T_10_addr] <= _T_fu_op__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_op1__T_10_en & _T_op1__T_10_mask) begin
      _T_op1[_T_op1__T_10_addr] <= _T_op1__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_id__T_10_en & _T_wb_id__T_10_mask) begin
      _T_wb_id[_T_wb_id__T_10_addr] <= _T_wb_id__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_pc__T_10_en & _T_wb_pc__T_10_mask) begin
      _T_wb_pc[_T_wb_pc__T_10_addr] <= _T_wb_pc__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_op__T_10_en & _T_wb_instr_op__T_10_mask) begin
      _T_wb_instr_op[_T_wb_instr_op__T_10_addr] <= _T_wb_instr_op__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_rs_idx__T_10_en & _T_wb_instr_rs_idx__T_10_mask) begin
      _T_wb_instr_rs_idx[_T_wb_instr_rs_idx__T_10_addr] <= _T_wb_instr_rs_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_rt_idx__T_10_en & _T_wb_instr_rt_idx__T_10_mask) begin
      _T_wb_instr_rt_idx[_T_wb_instr_rt_idx__T_10_addr] <= _T_wb_instr_rt_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_rd_idx__T_10_en & _T_wb_instr_rd_idx__T_10_mask) begin
      _T_wb_instr_rd_idx[_T_wb_instr_rd_idx__T_10_addr] <= _T_wb_instr_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_shamt__T_10_en & _T_wb_instr_shamt__T_10_mask) begin
      _T_wb_instr_shamt[_T_wb_instr_shamt__T_10_addr] <= _T_wb_instr_shamt__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_instr_func__T_10_en & _T_wb_instr_func__T_10_mask) begin
      _T_wb_instr_func[_T_wb_instr_func__T_10_addr] <= _T_wb_instr_func__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_rd_idx__T_10_en & _T_wb_rd_idx__T_10_mask) begin
      _T_wb_rd_idx[_T_wb_rd_idx__T_10_addr] <= _T_wb_rd_idx__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_ip7__T_10_en & _T_wb_ip7__T_10_mask) begin
      _T_wb_ip7[_T_wb_ip7__T_10_addr] <= _T_wb_ip7__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_is_ds__T_10_en & _T_wb_is_ds__T_10_mask) begin
      _T_wb_is_ds[_T_wb_is_ds__T_10_addr] <= _T_wb_is_ds__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_is_br__T_10_en & _T_wb_is_br__T_10_mask) begin
      _T_wb_is_br[_T_wb_is_br__T_10_addr] <= _T_wb_is_br__T_10_data; // @[Decoupled.scala 218:24]
    end
    if(_T_wb_npc__T_10_en & _T_wb_npc__T_10_mask) begin
      _T_wb_npc[_T_wb_npc__T_10_addr] <= _T_wb_npc__T_10_data; // @[Decoupled.scala 218:24]
    end
    if (reset) begin
      value <= 6'h0;
    end else if (_T_6) begin
      if (wrap) begin
        value <= 6'h0;
      end else begin
        value <= _T_12;
      end
    end
    if (reset) begin
      value_1 <= 6'h0;
    end else if (_T_8) begin
      if (wrap_1) begin
        value_1 <= 6'h0;
      end else begin
        value_1 <= _T_14;
      end
    end
    if (reset) begin
      _T_1 <= 1'h0;
    end else if (_T_15) begin
      _T_1 <= _T_6;
    end
  end
endmodule
module MDU_Divider(
  input         clock,
  input         reset,
  input         io_fu_in_valid,
  input  [5:0]  io_fu_in_bits_id,
  input  [4:0]  io_fu_in_bits_fu_op,
  input  [31:0] io_fu_in_bits_op1,
  input  [31:0] io_fu_in_bits_op2,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_ip7,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  output        io_fu_out_valid,
  output [5:0]  io_fu_out_bits_id,
  output [31:0] io_fu_out_bits_hi,
  output [31:0] io_fu_out_bits_lo,
  output [31:0] io_fu_out_bits_op1,
  output [4:0]  io_fu_out_bits_fu_op,
  output [7:0]  io_fu_out_bits_wb_id,
  output [31:0] io_fu_out_bits_wb_pc,
  output [5:0]  io_fu_out_bits_wb_instr_op,
  output [4:0]  io_fu_out_bits_wb_instr_rs_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rt_idx,
  output [4:0]  io_fu_out_bits_wb_instr_rd_idx,
  output [4:0]  io_fu_out_bits_wb_instr_shamt,
  output [5:0]  io_fu_out_bits_wb_instr_func,
  output [4:0]  io_fu_out_bits_wb_rd_idx,
  output        io_fu_out_bits_wb_ip7,
  output        io_fu_out_bits_wb_is_ds,
  output        io_fu_out_bits_wb_is_br,
  output [31:0] io_fu_out_bits_wb_npc,
  output        io_divider_data_dividend_tvalid,
  output        io_divider_data_divisor_tvalid,
  input         io_divider_data_dout_tvalid,
  output [39:0] io_divider_data_dividend_tdata,
  output [39:0] io_divider_data_divisor_tdata,
  input  [79:0] io_divider_data_dout_tdata
);
  wire  queue_clock; // @[mdu.scala 92:21]
  wire  queue_reset; // @[mdu.scala 92:21]
  wire  queue_io_enq_ready; // @[mdu.scala 92:21]
  wire  queue_io_enq_valid; // @[mdu.scala 92:21]
  wire [5:0] queue_io_enq_bits_id; // @[mdu.scala 92:21]
  wire [4:0] queue_io_enq_bits_fu_op; // @[mdu.scala 92:21]
  wire [31:0] queue_io_enq_bits_op1; // @[mdu.scala 92:21]
  wire [7:0] queue_io_enq_bits_wb_id; // @[mdu.scala 92:21]
  wire [31:0] queue_io_enq_bits_wb_pc; // @[mdu.scala 92:21]
  wire [5:0] queue_io_enq_bits_wb_instr_op; // @[mdu.scala 92:21]
  wire [4:0] queue_io_enq_bits_wb_instr_rs_idx; // @[mdu.scala 92:21]
  wire [4:0] queue_io_enq_bits_wb_instr_rt_idx; // @[mdu.scala 92:21]
  wire [4:0] queue_io_enq_bits_wb_instr_rd_idx; // @[mdu.scala 92:21]
  wire [4:0] queue_io_enq_bits_wb_instr_shamt; // @[mdu.scala 92:21]
  wire [5:0] queue_io_enq_bits_wb_instr_func; // @[mdu.scala 92:21]
  wire [4:0] queue_io_enq_bits_wb_rd_idx; // @[mdu.scala 92:21]
  wire  queue_io_enq_bits_wb_ip7; // @[mdu.scala 92:21]
  wire  queue_io_enq_bits_wb_is_ds; // @[mdu.scala 92:21]
  wire  queue_io_enq_bits_wb_is_br; // @[mdu.scala 92:21]
  wire [31:0] queue_io_enq_bits_wb_npc; // @[mdu.scala 92:21]
  wire  queue_io_deq_ready; // @[mdu.scala 92:21]
  wire  queue_io_deq_valid; // @[mdu.scala 92:21]
  wire [5:0] queue_io_deq_bits_id; // @[mdu.scala 92:21]
  wire [4:0] queue_io_deq_bits_fu_op; // @[mdu.scala 92:21]
  wire [31:0] queue_io_deq_bits_op1; // @[mdu.scala 92:21]
  wire [7:0] queue_io_deq_bits_wb_id; // @[mdu.scala 92:21]
  wire [31:0] queue_io_deq_bits_wb_pc; // @[mdu.scala 92:21]
  wire [5:0] queue_io_deq_bits_wb_instr_op; // @[mdu.scala 92:21]
  wire [4:0] queue_io_deq_bits_wb_instr_rs_idx; // @[mdu.scala 92:21]
  wire [4:0] queue_io_deq_bits_wb_instr_rt_idx; // @[mdu.scala 92:21]
  wire [4:0] queue_io_deq_bits_wb_instr_rd_idx; // @[mdu.scala 92:21]
  wire [4:0] queue_io_deq_bits_wb_instr_shamt; // @[mdu.scala 92:21]
  wire [5:0] queue_io_deq_bits_wb_instr_func; // @[mdu.scala 92:21]
  wire [4:0] queue_io_deq_bits_wb_rd_idx; // @[mdu.scala 92:21]
  wire  queue_io_deq_bits_wb_ip7; // @[mdu.scala 92:21]
  wire  queue_io_deq_bits_wb_is_ds; // @[mdu.scala 92:21]
  wire  queue_io_deq_bits_wb_is_br; // @[mdu.scala 92:21]
  wire [31:0] queue_io_deq_bits_wb_npc; // @[mdu.scala 92:21]
  wire  _T_3 = io_fu_in_bits_fu_op == 5'hf; // @[mdu.scala 105:47]
  wire [31:0] _T_5 = io_fu_in_bits_op1; // @[mdu.scala 106:17]
  wire [39:0] _T_6 = {{8{_T_5[31]}},_T_5}; // @[mdu.scala 106:30]
  wire [39:0] _T_7 = {{8'd0}, io_fu_in_bits_op1}; // @[mdu.scala 107:17 mdu.scala 107:17]
  wire [31:0] _T_11 = io_fu_in_bits_op2; // @[mdu.scala 109:17]
  wire [39:0] _T_12 = {{8{_T_11[31]}},_T_11}; // @[mdu.scala 109:30]
  wire [39:0] _T_13 = {{8'd0}, io_fu_in_bits_op2}; // @[mdu.scala 110:17 mdu.scala 110:17]
  Queue_1 queue ( // @[mdu.scala 92:21]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits_id(queue_io_enq_bits_id),
    .io_enq_bits_fu_op(queue_io_enq_bits_fu_op),
    .io_enq_bits_op1(queue_io_enq_bits_op1),
    .io_enq_bits_wb_id(queue_io_enq_bits_wb_id),
    .io_enq_bits_wb_pc(queue_io_enq_bits_wb_pc),
    .io_enq_bits_wb_instr_op(queue_io_enq_bits_wb_instr_op),
    .io_enq_bits_wb_instr_rs_idx(queue_io_enq_bits_wb_instr_rs_idx),
    .io_enq_bits_wb_instr_rt_idx(queue_io_enq_bits_wb_instr_rt_idx),
    .io_enq_bits_wb_instr_rd_idx(queue_io_enq_bits_wb_instr_rd_idx),
    .io_enq_bits_wb_instr_shamt(queue_io_enq_bits_wb_instr_shamt),
    .io_enq_bits_wb_instr_func(queue_io_enq_bits_wb_instr_func),
    .io_enq_bits_wb_rd_idx(queue_io_enq_bits_wb_rd_idx),
    .io_enq_bits_wb_ip7(queue_io_enq_bits_wb_ip7),
    .io_enq_bits_wb_is_ds(queue_io_enq_bits_wb_is_ds),
    .io_enq_bits_wb_is_br(queue_io_enq_bits_wb_is_br),
    .io_enq_bits_wb_npc(queue_io_enq_bits_wb_npc),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits_id(queue_io_deq_bits_id),
    .io_deq_bits_fu_op(queue_io_deq_bits_fu_op),
    .io_deq_bits_op1(queue_io_deq_bits_op1),
    .io_deq_bits_wb_id(queue_io_deq_bits_wb_id),
    .io_deq_bits_wb_pc(queue_io_deq_bits_wb_pc),
    .io_deq_bits_wb_instr_op(queue_io_deq_bits_wb_instr_op),
    .io_deq_bits_wb_instr_rs_idx(queue_io_deq_bits_wb_instr_rs_idx),
    .io_deq_bits_wb_instr_rt_idx(queue_io_deq_bits_wb_instr_rt_idx),
    .io_deq_bits_wb_instr_rd_idx(queue_io_deq_bits_wb_instr_rd_idx),
    .io_deq_bits_wb_instr_shamt(queue_io_deq_bits_wb_instr_shamt),
    .io_deq_bits_wb_instr_func(queue_io_deq_bits_wb_instr_func),
    .io_deq_bits_wb_rd_idx(queue_io_deq_bits_wb_rd_idx),
    .io_deq_bits_wb_ip7(queue_io_deq_bits_wb_ip7),
    .io_deq_bits_wb_is_ds(queue_io_deq_bits_wb_is_ds),
    .io_deq_bits_wb_is_br(queue_io_deq_bits_wb_is_br),
    .io_deq_bits_wb_npc(queue_io_deq_bits_wb_npc)
  );
  assign io_fu_out_valid = io_divider_data_dout_tvalid; // @[mdu.scala 113:19]
  assign io_fu_out_bits_id = queue_io_deq_bits_id; // @[mdu.scala 116:21]
  assign io_fu_out_bits_hi = io_divider_data_dout_tdata[31:0]; // @[mdu.scala 118:21]
  assign io_fu_out_bits_lo = io_divider_data_dout_tdata[71:40]; // @[mdu.scala 119:21]
  assign io_fu_out_bits_op1 = queue_io_deq_bits_op1; // @[mdu.scala 117:22]
  assign io_fu_out_bits_fu_op = queue_io_deq_bits_fu_op; // @[mdu.scala 115:24]
  assign io_fu_out_bits_wb_id = queue_io_deq_bits_wb_id; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_pc = queue_io_deq_bits_wb_pc; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_instr_op = queue_io_deq_bits_wb_instr_op; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_instr_rs_idx = queue_io_deq_bits_wb_instr_rs_idx; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_instr_rt_idx = queue_io_deq_bits_wb_instr_rt_idx; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_instr_rd_idx = queue_io_deq_bits_wb_instr_rd_idx; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_instr_shamt = queue_io_deq_bits_wb_instr_shamt; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_instr_func = queue_io_deq_bits_wb_instr_func; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_rd_idx = queue_io_deq_bits_wb_rd_idx; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_ip7 = queue_io_deq_bits_wb_ip7; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_is_ds = queue_io_deq_bits_wb_is_ds; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_is_br = queue_io_deq_bits_wb_is_br; // @[mdu.scala 114:21]
  assign io_fu_out_bits_wb_npc = queue_io_deq_bits_wb_npc; // @[mdu.scala 114:21]
  assign io_divider_data_dividend_tvalid = io_fu_in_valid; // @[mdu.scala 103:35]
  assign io_divider_data_divisor_tvalid = io_fu_in_valid; // @[mdu.scala 104:34]
  assign io_divider_data_dividend_tdata = _T_3 ? _T_6 : _T_7; // @[mdu.scala 105:34]
  assign io_divider_data_divisor_tdata = _T_3 ? _T_12 : _T_13; // @[mdu.scala 108:33]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = io_divider_data_dividend_tvalid & io_divider_data_divisor_tvalid; // @[mdu.scala 93:22]
  assign queue_io_enq_bits_id = io_fu_in_bits_id; // @[mdu.scala 94:24]
  assign queue_io_enq_bits_fu_op = io_fu_in_bits_fu_op; // @[mdu.scala 96:27]
  assign queue_io_enq_bits_op1 = io_fu_in_bits_op1; // @[mdu.scala 95:25]
  assign queue_io_enq_bits_wb_id = io_fu_in_bits_wb_id; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_pc = io_fu_in_bits_wb_pc; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_is_ds = io_fu_in_bits_wb_is_ds; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[mdu.scala 97:24]
  assign queue_io_enq_bits_wb_npc = io_fu_in_bits_wb_npc; // @[mdu.scala 97:24]
  assign queue_io_deq_ready = io_divider_data_dout_tvalid; // @[mdu.scala 98:22]
endmodule
module ROB(
  input         clock,
  input         reset,
  input         io_enq_0_valid,
  input  [5:0]  io_enq_0_bits_id,
  input  [31:0] io_enq_0_bits_data_hi,
  input  [31:0] io_enq_0_bits_data_lo,
  input  [31:0] io_enq_0_bits_data_op1,
  input  [4:0]  io_enq_0_bits_data_fu_op,
  input  [7:0]  io_enq_0_bits_data_wb_id,
  input  [31:0] io_enq_0_bits_data_wb_pc,
  input  [5:0]  io_enq_0_bits_data_wb_instr_op,
  input  [4:0]  io_enq_0_bits_data_wb_instr_rs_idx,
  input  [4:0]  io_enq_0_bits_data_wb_instr_rt_idx,
  input  [4:0]  io_enq_0_bits_data_wb_instr_rd_idx,
  input  [4:0]  io_enq_0_bits_data_wb_instr_shamt,
  input  [5:0]  io_enq_0_bits_data_wb_instr_func,
  input  [4:0]  io_enq_0_bits_data_wb_rd_idx,
  input         io_enq_0_bits_data_wb_ip7,
  input         io_enq_0_bits_data_wb_is_ds,
  input         io_enq_0_bits_data_wb_is_br,
  input  [31:0] io_enq_0_bits_data_wb_npc,
  input         io_enq_1_valid,
  input  [5:0]  io_enq_1_bits_id,
  input  [31:0] io_enq_1_bits_data_hi,
  input  [31:0] io_enq_1_bits_data_lo,
  input  [31:0] io_enq_1_bits_data_op1,
  input  [4:0]  io_enq_1_bits_data_fu_op,
  input  [7:0]  io_enq_1_bits_data_wb_id,
  input  [31:0] io_enq_1_bits_data_wb_pc,
  input  [5:0]  io_enq_1_bits_data_wb_instr_op,
  input  [4:0]  io_enq_1_bits_data_wb_instr_rs_idx,
  input  [4:0]  io_enq_1_bits_data_wb_instr_rt_idx,
  input  [4:0]  io_enq_1_bits_data_wb_instr_rd_idx,
  input  [4:0]  io_enq_1_bits_data_wb_instr_shamt,
  input  [5:0]  io_enq_1_bits_data_wb_instr_func,
  input  [4:0]  io_enq_1_bits_data_wb_rd_idx,
  input         io_enq_1_bits_data_wb_ip7,
  input         io_enq_1_bits_data_wb_is_ds,
  input         io_enq_1_bits_data_wb_is_br,
  input  [31:0] io_enq_1_bits_data_wb_npc,
  output        io_deq_valid,
  output [31:0] io_deq_bits_hi,
  output [31:0] io_deq_bits_lo,
  output [31:0] io_deq_bits_op1,
  output [4:0]  io_deq_bits_fu_op,
  output [7:0]  io_deq_bits_wb_id,
  output [31:0] io_deq_bits_wb_pc,
  output [5:0]  io_deq_bits_wb_instr_op,
  output [4:0]  io_deq_bits_wb_instr_rs_idx,
  output [4:0]  io_deq_bits_wb_instr_rt_idx,
  output [4:0]  io_deq_bits_wb_instr_rd_idx,
  output [4:0]  io_deq_bits_wb_instr_shamt,
  output [5:0]  io_deq_bits_wb_instr_func,
  output [4:0]  io_deq_bits_wb_rd_idx,
  output        io_deq_bits_wb_ip7,
  output        io_deq_bits_wb_is_ds,
  output        io_deq_bits_wb_is_br,
  output [31:0] io_deq_bits_wb_npc
);
  reg  queue_valid [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_0;
  wire  queue_valid_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid_q_head_r_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_3_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_3_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_3_en; // @[utils.scala 30:18]
  wire  queue_valid__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_4_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_4_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_4_en; // @[utils.scala 30:18]
  wire  queue_valid__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_5_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_5_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_5_en; // @[utils.scala 30:18]
  wire  queue_valid__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_6_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_6_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_6_en; // @[utils.scala 30:18]
  wire  queue_valid__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_7_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_7_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_7_en; // @[utils.scala 30:18]
  wire  queue_valid__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_8_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_8_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_8_en; // @[utils.scala 30:18]
  wire  queue_valid__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_9_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_9_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_9_en; // @[utils.scala 30:18]
  wire  queue_valid__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_10_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_10_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_10_en; // @[utils.scala 30:18]
  wire  queue_valid__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_11_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_11_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_11_en; // @[utils.scala 30:18]
  wire  queue_valid__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_12_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_12_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_12_en; // @[utils.scala 30:18]
  wire  queue_valid__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_13_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_13_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_13_en; // @[utils.scala 30:18]
  wire  queue_valid__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_14_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_14_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_14_en; // @[utils.scala 30:18]
  wire  queue_valid__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_15_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_15_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_15_en; // @[utils.scala 30:18]
  wire  queue_valid__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_16_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_16_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_16_en; // @[utils.scala 30:18]
  wire  queue_valid__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_17_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_17_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_17_en; // @[utils.scala 30:18]
  wire  queue_valid__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_18_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_18_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_18_en; // @[utils.scala 30:18]
  wire  queue_valid__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_19_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_19_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_19_en; // @[utils.scala 30:18]
  wire  queue_valid__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_20_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_20_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_20_en; // @[utils.scala 30:18]
  wire  queue_valid__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_21_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_21_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_21_en; // @[utils.scala 30:18]
  wire  queue_valid__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_22_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_22_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_22_en; // @[utils.scala 30:18]
  wire  queue_valid__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_23_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_23_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_23_en; // @[utils.scala 30:18]
  wire  queue_valid__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_24_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_24_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_24_en; // @[utils.scala 30:18]
  wire  queue_valid__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_25_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_25_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_25_en; // @[utils.scala 30:18]
  wire  queue_valid__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_26_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_26_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_26_en; // @[utils.scala 30:18]
  wire  queue_valid__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_27_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_27_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_27_en; // @[utils.scala 30:18]
  wire  queue_valid__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_28_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_28_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_28_en; // @[utils.scala 30:18]
  wire  queue_valid__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_29_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_29_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_29_en; // @[utils.scala 30:18]
  wire  queue_valid__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_30_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_30_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_30_en; // @[utils.scala 30:18]
  wire  queue_valid__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_31_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_31_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_31_en; // @[utils.scala 30:18]
  wire  queue_valid__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_32_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_32_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_32_en; // @[utils.scala 30:18]
  wire  queue_valid__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_33_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_33_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_33_en; // @[utils.scala 30:18]
  wire  queue_valid__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_34_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_34_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_34_en; // @[utils.scala 30:18]
  wire  queue_valid__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_35_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_35_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_35_en; // @[utils.scala 30:18]
  wire  queue_valid__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_36_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_36_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_36_en; // @[utils.scala 30:18]
  wire  queue_valid__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_37_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_37_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_37_en; // @[utils.scala 30:18]
  wire  queue_valid__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_38_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_38_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_38_en; // @[utils.scala 30:18]
  wire  queue_valid__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_39_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_39_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_39_en; // @[utils.scala 30:18]
  wire  queue_valid__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_40_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_40_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_40_en; // @[utils.scala 30:18]
  wire  queue_valid__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_41_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_41_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_41_en; // @[utils.scala 30:18]
  wire  queue_valid__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_42_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_42_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_42_en; // @[utils.scala 30:18]
  wire  queue_valid__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_43_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_43_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_43_en; // @[utils.scala 30:18]
  wire  queue_valid__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_44_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_44_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_44_en; // @[utils.scala 30:18]
  wire  queue_valid__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_45_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_45_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_45_en; // @[utils.scala 30:18]
  wire  queue_valid__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_46_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_46_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_46_en; // @[utils.scala 30:18]
  wire  queue_valid__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_47_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_47_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_47_en; // @[utils.scala 30:18]
  wire  queue_valid__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_48_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_48_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_48_en; // @[utils.scala 30:18]
  wire  queue_valid__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_49_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_49_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_49_en; // @[utils.scala 30:18]
  wire  queue_valid__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_50_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_50_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_50_en; // @[utils.scala 30:18]
  wire  queue_valid__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_51_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_51_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_51_en; // @[utils.scala 30:18]
  wire  queue_valid__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_52_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_52_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_52_en; // @[utils.scala 30:18]
  wire  queue_valid__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_53_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_53_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_53_en; // @[utils.scala 30:18]
  wire  queue_valid__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_54_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_54_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_54_en; // @[utils.scala 30:18]
  wire  queue_valid__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_55_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_55_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_55_en; // @[utils.scala 30:18]
  wire  queue_valid__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_56_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_56_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_56_en; // @[utils.scala 30:18]
  wire  queue_valid__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_57_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_57_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_57_en; // @[utils.scala 30:18]
  wire  queue_valid__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_58_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_58_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_58_en; // @[utils.scala 30:18]
  wire  queue_valid__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_59_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_59_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_59_en; // @[utils.scala 30:18]
  wire  queue_valid__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_60_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_60_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_60_en; // @[utils.scala 30:18]
  wire  queue_valid__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_61_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_61_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_61_en; // @[utils.scala 30:18]
  wire  queue_valid__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_62_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_62_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_62_en; // @[utils.scala 30:18]
  wire  queue_valid__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_63_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_63_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_63_en; // @[utils.scala 30:18]
  wire  queue_valid__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_64_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_64_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_64_en; // @[utils.scala 30:18]
  wire  queue_valid__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_65_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_65_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_65_en; // @[utils.scala 30:18]
  wire  queue_valid__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_66_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_66_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_66_en; // @[utils.scala 30:18]
  wire  queue_valid__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_67_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_67_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_67_en; // @[utils.scala 30:18]
  wire  queue_valid__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_68_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_68_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_68_en; // @[utils.scala 30:18]
  wire  queue_valid__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_70_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_70_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_70_en; // @[utils.scala 30:18]
  wire  queue_valid__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_71_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_71_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_71_en; // @[utils.scala 30:18]
  wire  queue_valid__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_72_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_72_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_72_en; // @[utils.scala 30:18]
  wire  queue_valid__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_73_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_73_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_73_en; // @[utils.scala 30:18]
  wire  queue_valid__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_74_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_74_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_74_en; // @[utils.scala 30:18]
  wire  queue_valid__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_75_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_75_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_75_en; // @[utils.scala 30:18]
  wire  queue_valid__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_76_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_76_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_76_en; // @[utils.scala 30:18]
  wire  queue_valid__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_77_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_77_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_77_en; // @[utils.scala 30:18]
  wire  queue_valid__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_78_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_78_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_78_en; // @[utils.scala 30:18]
  wire  queue_valid__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_79_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_79_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_79_en; // @[utils.scala 30:18]
  wire  queue_valid__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_80_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_80_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_80_en; // @[utils.scala 30:18]
  wire  queue_valid__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_81_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_81_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_81_en; // @[utils.scala 30:18]
  wire  queue_valid__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_82_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_82_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_82_en; // @[utils.scala 30:18]
  wire  queue_valid__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_83_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_83_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_83_en; // @[utils.scala 30:18]
  wire  queue_valid__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_84_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_84_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_84_en; // @[utils.scala 30:18]
  wire  queue_valid__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_85_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_85_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_85_en; // @[utils.scala 30:18]
  wire  queue_valid__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_86_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_86_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_86_en; // @[utils.scala 30:18]
  wire  queue_valid__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_87_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_87_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_87_en; // @[utils.scala 30:18]
  wire  queue_valid__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_88_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_88_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_88_en; // @[utils.scala 30:18]
  wire  queue_valid__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_89_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_89_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_89_en; // @[utils.scala 30:18]
  wire  queue_valid__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_90_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_90_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_90_en; // @[utils.scala 30:18]
  wire  queue_valid__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_91_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_91_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_91_en; // @[utils.scala 30:18]
  wire  queue_valid__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_92_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_92_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_92_en; // @[utils.scala 30:18]
  wire  queue_valid__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_93_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_93_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_93_en; // @[utils.scala 30:18]
  wire  queue_valid__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_94_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_94_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_94_en; // @[utils.scala 30:18]
  wire  queue_valid__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_95_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_95_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_95_en; // @[utils.scala 30:18]
  wire  queue_valid__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_96_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_96_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_96_en; // @[utils.scala 30:18]
  wire  queue_valid__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_97_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_97_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_97_en; // @[utils.scala 30:18]
  wire  queue_valid__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_98_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_98_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_98_en; // @[utils.scala 30:18]
  wire  queue_valid__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_99_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_99_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_99_en; // @[utils.scala 30:18]
  wire  queue_valid__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_100_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_100_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_100_en; // @[utils.scala 30:18]
  wire  queue_valid__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_101_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_101_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_101_en; // @[utils.scala 30:18]
  wire  queue_valid__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_102_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_102_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_102_en; // @[utils.scala 30:18]
  wire  queue_valid__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_103_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_103_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_103_en; // @[utils.scala 30:18]
  wire  queue_valid__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_104_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_104_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_104_en; // @[utils.scala 30:18]
  wire  queue_valid__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_105_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_105_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_105_en; // @[utils.scala 30:18]
  wire  queue_valid__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_106_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_106_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_106_en; // @[utils.scala 30:18]
  wire  queue_valid__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_107_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_107_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_107_en; // @[utils.scala 30:18]
  wire  queue_valid__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_108_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_108_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_108_en; // @[utils.scala 30:18]
  wire  queue_valid__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_109_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_109_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_109_en; // @[utils.scala 30:18]
  wire  queue_valid__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_110_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_110_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_110_en; // @[utils.scala 30:18]
  wire  queue_valid__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_111_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_111_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_111_en; // @[utils.scala 30:18]
  wire  queue_valid__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_112_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_112_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_112_en; // @[utils.scala 30:18]
  wire  queue_valid__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_113_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_113_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_113_en; // @[utils.scala 30:18]
  wire  queue_valid__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_114_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_114_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_114_en; // @[utils.scala 30:18]
  wire  queue_valid__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_115_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_115_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_115_en; // @[utils.scala 30:18]
  wire  queue_valid__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_116_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_116_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_116_en; // @[utils.scala 30:18]
  wire  queue_valid__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_117_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_117_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_117_en; // @[utils.scala 30:18]
  wire  queue_valid__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_118_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_118_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_118_en; // @[utils.scala 30:18]
  wire  queue_valid__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_119_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_119_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_119_en; // @[utils.scala 30:18]
  wire  queue_valid__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_120_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_120_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_120_en; // @[utils.scala 30:18]
  wire  queue_valid__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_121_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_121_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_121_en; // @[utils.scala 30:18]
  wire  queue_valid__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_122_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_122_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_122_en; // @[utils.scala 30:18]
  wire  queue_valid__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_123_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_123_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_123_en; // @[utils.scala 30:18]
  wire  queue_valid__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_124_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_124_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_124_en; // @[utils.scala 30:18]
  wire  queue_valid__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_125_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_125_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_125_en; // @[utils.scala 30:18]
  wire  queue_valid__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_126_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_126_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_126_en; // @[utils.scala 30:18]
  wire  queue_valid__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_127_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_127_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_127_en; // @[utils.scala 30:18]
  wire  queue_valid__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_128_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_128_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_128_en; // @[utils.scala 30:18]
  wire  queue_valid__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_129_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_129_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_129_en; // @[utils.scala 30:18]
  wire  queue_valid__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_130_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_130_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_130_en; // @[utils.scala 30:18]
  wire  queue_valid__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_131_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_131_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_131_en; // @[utils.scala 30:18]
  wire  queue_valid__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_132_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_132_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_132_en; // @[utils.scala 30:18]
  wire  queue_valid__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid__T_133_addr; // @[utils.scala 30:18]
  wire  queue_valid__T_133_mask; // @[utils.scala 30:18]
  wire  queue_valid__T_133_en; // @[utils.scala 30:18]
  wire  queue_valid_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_valid_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_valid_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_valid_q_head_w_en; // @[utils.scala 30:18]
  reg [31:0] queue_bits_hi [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_1;
  wire [31:0] queue_bits_hi_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi_q_head_r_addr; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_3_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_4_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_5_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_6_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_7_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_8_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_9_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_10_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_11_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_12_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_13_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_14_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_15_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_16_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_17_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_18_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_19_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_20_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_21_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_22_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_23_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_24_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_25_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_26_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_27_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_28_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_29_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_30_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_31_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_32_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_33_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_34_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_35_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_36_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_37_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_38_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_39_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_40_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_41_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_42_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_43_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_44_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_45_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_46_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_47_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_48_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_49_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_50_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_51_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_52_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_53_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_54_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_55_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_56_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_57_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_58_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_59_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_60_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_61_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_62_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_63_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_64_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_65_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_66_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_67_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_68_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_70_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_71_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_72_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_73_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_74_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_75_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_76_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_77_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_78_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_79_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_80_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_81_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_82_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_83_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_84_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_85_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_86_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_87_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_88_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_89_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_90_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_91_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_92_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_93_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_94_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_95_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_96_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_97_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_98_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_99_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_100_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_101_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_102_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_103_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_104_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_105_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_106_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_107_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_108_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_109_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_110_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_111_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_112_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_113_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_114_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_115_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_116_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_117_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_118_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_119_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_120_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_121_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_122_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_123_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_124_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_125_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_126_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_127_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_128_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_129_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_130_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_131_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_132_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi__T_133_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_hi_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_hi_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_hi_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_hi_q_head_w_en; // @[utils.scala 30:18]
  reg [31:0] queue_bits_lo [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_2;
  wire [31:0] queue_bits_lo_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo_q_head_r_addr; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_3_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_4_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_5_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_6_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_7_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_8_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_9_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_10_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_11_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_12_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_13_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_14_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_15_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_16_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_17_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_18_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_19_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_20_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_21_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_22_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_23_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_24_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_25_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_26_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_27_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_28_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_29_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_30_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_31_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_32_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_33_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_34_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_35_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_36_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_37_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_38_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_39_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_40_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_41_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_42_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_43_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_44_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_45_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_46_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_47_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_48_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_49_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_50_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_51_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_52_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_53_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_54_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_55_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_56_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_57_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_58_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_59_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_60_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_61_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_62_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_63_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_64_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_65_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_66_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_67_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_68_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_70_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_71_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_72_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_73_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_74_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_75_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_76_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_77_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_78_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_79_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_80_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_81_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_82_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_83_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_84_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_85_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_86_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_87_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_88_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_89_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_90_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_91_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_92_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_93_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_94_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_95_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_96_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_97_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_98_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_99_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_100_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_101_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_102_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_103_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_104_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_105_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_106_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_107_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_108_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_109_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_110_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_111_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_112_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_113_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_114_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_115_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_116_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_117_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_118_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_119_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_120_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_121_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_122_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_123_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_124_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_125_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_126_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_127_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_128_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_129_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_130_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_131_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_132_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo__T_133_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_lo_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_lo_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_lo_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_lo_q_head_w_en; // @[utils.scala 30:18]
  reg [31:0] queue_bits_op1 [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_3;
  wire [31:0] queue_bits_op1_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1_q_head_r_addr; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_3_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_4_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_5_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_6_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_7_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_8_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_9_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_10_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_11_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_12_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_13_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_14_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_15_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_16_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_17_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_18_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_19_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_20_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_21_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_22_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_23_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_24_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_25_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_26_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_27_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_28_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_29_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_30_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_31_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_32_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_33_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_34_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_35_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_36_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_37_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_38_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_39_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_40_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_41_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_42_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_43_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_44_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_45_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_46_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_47_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_48_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_49_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_50_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_51_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_52_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_53_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_54_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_55_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_56_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_57_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_58_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_59_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_60_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_61_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_62_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_63_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_64_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_65_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_66_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_67_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_68_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_70_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_71_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_72_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_73_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_74_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_75_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_76_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_77_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_78_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_79_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_80_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_81_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_82_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_83_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_84_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_85_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_86_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_87_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_88_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_89_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_90_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_91_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_92_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_93_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_94_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_95_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_96_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_97_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_98_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_99_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_100_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_101_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_102_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_103_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_104_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_105_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_106_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_107_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_108_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_109_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_110_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_111_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_112_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_113_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_114_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_115_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_116_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_117_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_118_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_119_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_120_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_121_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_122_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_123_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_124_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_125_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_126_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_127_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_128_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_129_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_130_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_131_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_132_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1__T_133_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_op1_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_op1_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_op1_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_op1_q_head_w_en; // @[utils.scala 30:18]
  reg [4:0] queue_bits_fu_op [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_4;
  wire [4:0] queue_bits_fu_op_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op_q_head_r_addr; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_3_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_4_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_5_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_6_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_7_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_8_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_9_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_10_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_11_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_12_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_13_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_14_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_15_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_16_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_17_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_18_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_19_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_20_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_21_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_22_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_23_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_24_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_25_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_26_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_27_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_28_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_29_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_30_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_31_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_32_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_33_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_34_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_35_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_36_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_37_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_38_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_39_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_40_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_41_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_42_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_43_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_44_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_45_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_46_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_47_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_48_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_49_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_50_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_51_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_52_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_53_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_54_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_55_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_56_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_57_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_58_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_59_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_60_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_61_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_62_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_63_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_64_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_65_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_66_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_67_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_68_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_70_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_71_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_72_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_73_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_74_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_75_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_76_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_77_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_78_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_79_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_80_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_81_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_82_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_83_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_84_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_85_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_86_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_87_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_88_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_89_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_90_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_91_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_92_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_93_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_94_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_95_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_96_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_97_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_98_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_99_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_100_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_101_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_102_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_103_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_104_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_105_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_106_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_107_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_108_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_109_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_110_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_111_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_112_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_113_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_114_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_115_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_116_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_117_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_118_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_119_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_120_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_121_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_122_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_123_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_124_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_125_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_126_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_127_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_128_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_129_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_130_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_131_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_132_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op__T_133_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_fu_op_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_fu_op_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_fu_op_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_fu_op_q_head_w_en; // @[utils.scala 30:18]
  reg [7:0] queue_bits_wb_id [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_5;
  wire [7:0] queue_bits_wb_id_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id_q_head_r_addr; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_3_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_4_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_5_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_6_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_7_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_8_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_9_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_10_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_11_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_12_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_13_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_14_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_15_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_16_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_17_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_18_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_19_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_20_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_21_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_22_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_23_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_24_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_25_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_26_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_27_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_28_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_29_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_30_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_31_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_32_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_33_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_34_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_35_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_36_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_37_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_38_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_39_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_40_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_41_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_42_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_43_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_44_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_45_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_46_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_47_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_48_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_49_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_50_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_51_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_52_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_53_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_54_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_55_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_56_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_57_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_58_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_59_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_60_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_61_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_62_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_63_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_64_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_65_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_66_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_67_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_68_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_70_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_71_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_72_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_73_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_74_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_75_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_76_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_77_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_78_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_79_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_80_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_81_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_82_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_83_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_84_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_85_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_86_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_87_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_88_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_89_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_90_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_91_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_92_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_93_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_94_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_95_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_96_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_97_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_98_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_99_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_100_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_101_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_102_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_103_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_104_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_105_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_106_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_107_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_108_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_109_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_110_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_111_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_112_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_113_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_114_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_115_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_116_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_117_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_118_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_119_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_120_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_121_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_122_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_123_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_124_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_125_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_126_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_127_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_128_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_129_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_130_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_131_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_132_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id__T_133_en; // @[utils.scala 30:18]
  wire [7:0] queue_bits_wb_id_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_id_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_id_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_id_q_head_w_en; // @[utils.scala 30:18]
  reg [31:0] queue_bits_wb_pc [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_6;
  wire [31:0] queue_bits_wb_pc_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc_q_head_r_addr; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_3_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_4_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_5_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_6_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_7_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_8_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_9_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_10_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_11_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_12_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_13_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_14_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_15_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_16_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_17_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_18_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_19_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_20_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_21_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_22_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_23_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_24_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_25_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_26_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_27_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_28_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_29_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_30_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_31_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_32_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_33_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_34_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_35_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_36_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_37_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_38_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_39_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_40_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_41_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_42_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_43_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_44_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_45_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_46_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_47_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_48_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_49_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_50_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_51_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_52_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_53_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_54_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_55_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_56_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_57_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_58_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_59_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_60_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_61_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_62_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_63_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_64_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_65_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_66_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_67_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_68_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_70_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_71_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_72_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_73_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_74_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_75_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_76_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_77_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_78_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_79_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_80_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_81_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_82_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_83_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_84_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_85_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_86_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_87_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_88_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_89_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_90_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_91_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_92_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_93_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_94_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_95_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_96_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_97_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_98_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_99_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_100_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_101_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_102_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_103_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_104_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_105_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_106_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_107_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_108_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_109_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_110_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_111_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_112_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_113_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_114_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_115_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_116_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_117_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_118_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_119_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_120_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_121_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_122_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_123_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_124_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_125_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_126_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_127_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_128_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_129_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_130_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_131_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_132_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc__T_133_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_pc_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_pc_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_pc_q_head_w_en; // @[utils.scala 30:18]
  reg [5:0] queue_bits_wb_instr_op [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_7;
  wire [5:0] queue_bits_wb_instr_op_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op_q_head_r_addr; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_3_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_4_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_5_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_6_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_7_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_8_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_9_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_10_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_11_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_12_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_13_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_14_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_15_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_16_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_17_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_18_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_19_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_20_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_21_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_22_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_23_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_24_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_25_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_26_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_27_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_28_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_29_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_30_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_31_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_32_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_33_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_34_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_35_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_36_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_37_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_38_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_39_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_40_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_41_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_42_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_43_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_44_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_45_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_46_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_47_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_48_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_49_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_50_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_51_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_52_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_53_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_54_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_55_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_56_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_57_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_58_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_59_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_60_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_61_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_62_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_63_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_64_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_65_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_66_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_67_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_68_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_70_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_71_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_72_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_73_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_74_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_75_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_76_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_77_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_78_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_79_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_80_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_81_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_82_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_83_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_84_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_85_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_86_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_87_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_88_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_89_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_90_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_91_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_92_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_93_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_94_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_95_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_96_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_97_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_98_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_99_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_100_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_101_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_102_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_103_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_104_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_105_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_106_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_107_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_108_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_109_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_110_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_111_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_112_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_113_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_114_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_115_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_116_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_117_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_118_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_119_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_120_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_121_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_122_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_123_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_124_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_125_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_126_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_127_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_128_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_129_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_130_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_131_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_132_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op__T_133_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_op_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_op_q_head_w_en; // @[utils.scala 30:18]
  reg [4:0] queue_bits_wb_instr_rs_idx [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_8;
  wire [4:0] queue_bits_wb_instr_rs_idx_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx_q_head_r_addr; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_3_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_4_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_5_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_6_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_7_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_8_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_9_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_10_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_11_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_12_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_13_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_14_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_15_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_16_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_17_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_18_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_19_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_20_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_21_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_22_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_23_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_24_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_25_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_26_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_27_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_28_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_29_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_30_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_31_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_32_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_33_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_34_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_35_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_36_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_37_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_38_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_39_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_40_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_41_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_42_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_43_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_44_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_45_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_46_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_47_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_48_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_49_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_50_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_51_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_52_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_53_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_54_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_55_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_56_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_57_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_58_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_59_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_60_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_61_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_62_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_63_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_64_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_65_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_66_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_67_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_68_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_70_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_71_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_72_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_73_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_74_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_75_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_76_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_77_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_78_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_79_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_80_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_81_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_82_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_83_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_84_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_85_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_86_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_87_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_88_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_89_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_90_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_91_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_92_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_93_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_94_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_95_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_96_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_97_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_98_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_99_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_100_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_101_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_102_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_103_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_104_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_105_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_106_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_107_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_108_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_109_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_110_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_111_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_112_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_113_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_114_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_115_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_116_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_117_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_118_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_119_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_120_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_121_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_122_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_123_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_124_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_125_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_126_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_127_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_128_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_129_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_130_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_131_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_132_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx__T_133_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rs_idx_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rs_idx_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rs_idx_q_head_w_en; // @[utils.scala 30:18]
  reg [4:0] queue_bits_wb_instr_rt_idx [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_9;
  wire [4:0] queue_bits_wb_instr_rt_idx_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx_q_head_r_addr; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_3_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_4_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_5_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_6_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_7_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_8_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_9_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_10_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_11_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_12_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_13_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_14_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_15_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_16_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_17_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_18_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_19_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_20_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_21_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_22_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_23_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_24_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_25_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_26_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_27_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_28_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_29_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_30_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_31_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_32_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_33_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_34_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_35_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_36_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_37_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_38_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_39_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_40_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_41_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_42_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_43_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_44_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_45_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_46_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_47_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_48_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_49_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_50_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_51_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_52_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_53_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_54_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_55_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_56_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_57_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_58_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_59_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_60_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_61_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_62_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_63_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_64_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_65_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_66_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_67_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_68_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_70_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_71_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_72_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_73_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_74_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_75_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_76_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_77_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_78_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_79_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_80_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_81_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_82_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_83_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_84_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_85_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_86_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_87_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_88_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_89_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_90_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_91_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_92_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_93_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_94_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_95_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_96_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_97_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_98_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_99_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_100_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_101_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_102_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_103_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_104_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_105_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_106_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_107_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_108_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_109_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_110_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_111_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_112_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_113_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_114_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_115_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_116_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_117_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_118_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_119_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_120_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_121_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_122_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_123_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_124_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_125_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_126_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_127_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_128_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_129_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_130_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_131_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_132_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx__T_133_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rt_idx_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rt_idx_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rt_idx_q_head_w_en; // @[utils.scala 30:18]
  reg [4:0] queue_bits_wb_instr_rd_idx [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_10;
  wire [4:0] queue_bits_wb_instr_rd_idx_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx_q_head_r_addr; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_3_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_4_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_5_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_6_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_7_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_8_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_9_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_10_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_11_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_12_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_13_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_14_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_15_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_16_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_17_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_18_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_19_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_20_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_21_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_22_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_23_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_24_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_25_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_26_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_27_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_28_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_29_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_30_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_31_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_32_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_33_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_34_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_35_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_36_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_37_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_38_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_39_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_40_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_41_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_42_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_43_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_44_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_45_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_46_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_47_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_48_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_49_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_50_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_51_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_52_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_53_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_54_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_55_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_56_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_57_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_58_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_59_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_60_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_61_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_62_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_63_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_64_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_65_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_66_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_67_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_68_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_70_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_71_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_72_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_73_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_74_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_75_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_76_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_77_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_78_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_79_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_80_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_81_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_82_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_83_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_84_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_85_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_86_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_87_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_88_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_89_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_90_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_91_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_92_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_93_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_94_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_95_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_96_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_97_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_98_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_99_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_100_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_101_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_102_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_103_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_104_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_105_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_106_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_107_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_108_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_109_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_110_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_111_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_112_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_113_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_114_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_115_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_116_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_117_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_118_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_119_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_120_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_121_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_122_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_123_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_124_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_125_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_126_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_127_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_128_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_129_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_130_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_131_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_132_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx__T_133_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_rd_idx_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_rd_idx_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_rd_idx_q_head_w_en; // @[utils.scala 30:18]
  reg [4:0] queue_bits_wb_instr_shamt [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_11;
  wire [4:0] queue_bits_wb_instr_shamt_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt_q_head_r_addr; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_3_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_4_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_5_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_6_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_7_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_8_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_9_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_10_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_11_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_12_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_13_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_14_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_15_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_16_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_17_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_18_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_19_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_20_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_21_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_22_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_23_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_24_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_25_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_26_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_27_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_28_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_29_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_30_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_31_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_32_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_33_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_34_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_35_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_36_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_37_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_38_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_39_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_40_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_41_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_42_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_43_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_44_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_45_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_46_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_47_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_48_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_49_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_50_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_51_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_52_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_53_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_54_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_55_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_56_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_57_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_58_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_59_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_60_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_61_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_62_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_63_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_64_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_65_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_66_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_67_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_68_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_70_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_71_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_72_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_73_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_74_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_75_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_76_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_77_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_78_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_79_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_80_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_81_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_82_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_83_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_84_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_85_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_86_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_87_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_88_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_89_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_90_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_91_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_92_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_93_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_94_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_95_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_96_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_97_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_98_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_99_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_100_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_101_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_102_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_103_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_104_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_105_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_106_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_107_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_108_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_109_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_110_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_111_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_112_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_113_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_114_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_115_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_116_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_117_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_118_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_119_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_120_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_121_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_122_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_123_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_124_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_125_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_126_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_127_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_128_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_129_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_130_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_131_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_132_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt__T_133_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_instr_shamt_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_shamt_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_shamt_q_head_w_en; // @[utils.scala 30:18]
  reg [5:0] queue_bits_wb_instr_func [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_12;
  wire [5:0] queue_bits_wb_instr_func_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func_q_head_r_addr; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_3_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_4_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_5_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_6_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_7_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_8_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_9_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_10_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_11_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_12_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_13_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_14_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_15_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_16_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_17_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_18_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_19_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_20_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_21_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_22_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_23_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_24_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_25_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_26_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_27_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_28_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_29_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_30_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_31_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_32_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_33_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_34_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_35_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_36_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_37_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_38_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_39_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_40_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_41_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_42_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_43_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_44_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_45_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_46_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_47_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_48_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_49_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_50_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_51_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_52_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_53_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_54_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_55_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_56_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_57_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_58_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_59_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_60_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_61_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_62_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_63_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_64_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_65_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_66_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_67_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_68_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_70_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_71_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_72_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_73_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_74_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_75_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_76_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_77_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_78_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_79_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_80_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_81_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_82_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_83_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_84_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_85_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_86_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_87_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_88_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_89_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_90_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_91_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_92_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_93_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_94_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_95_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_96_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_97_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_98_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_99_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_100_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_101_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_102_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_103_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_104_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_105_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_106_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_107_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_108_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_109_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_110_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_111_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_112_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_113_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_114_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_115_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_116_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_117_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_118_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_119_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_120_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_121_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_122_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_123_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_124_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_125_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_126_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_127_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_128_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_129_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_130_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_131_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_132_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func__T_133_en; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_instr_func_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_instr_func_q_head_w_en; // @[utils.scala 30:18]
  reg [4:0] queue_bits_wb_rd_idx [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_13;
  wire [4:0] queue_bits_wb_rd_idx_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx_q_head_r_addr; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_3_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_4_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_5_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_6_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_7_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_8_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_9_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_10_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_11_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_12_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_13_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_14_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_15_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_16_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_17_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_18_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_19_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_20_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_21_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_22_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_23_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_24_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_25_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_26_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_27_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_28_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_29_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_30_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_31_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_32_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_33_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_34_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_35_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_36_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_37_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_38_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_39_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_40_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_41_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_42_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_43_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_44_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_45_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_46_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_47_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_48_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_49_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_50_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_51_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_52_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_53_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_54_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_55_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_56_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_57_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_58_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_59_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_60_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_61_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_62_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_63_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_64_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_65_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_66_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_67_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_68_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_70_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_71_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_72_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_73_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_74_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_75_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_76_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_77_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_78_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_79_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_80_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_81_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_82_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_83_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_84_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_85_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_86_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_87_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_88_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_89_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_90_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_91_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_92_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_93_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_94_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_95_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_96_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_97_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_98_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_99_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_100_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_101_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_102_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_103_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_104_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_105_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_106_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_107_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_108_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_109_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_110_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_111_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_112_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_113_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_114_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_115_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_116_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_117_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_118_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_119_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_120_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_121_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_122_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_123_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_124_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_125_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_126_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_127_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_128_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_129_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_130_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_131_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_132_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx__T_133_en; // @[utils.scala 30:18]
  wire [4:0] queue_bits_wb_rd_idx_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_rd_idx_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_rd_idx_q_head_w_en; // @[utils.scala 30:18]
  reg  queue_bits_wb_ip7 [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_14;
  wire  queue_bits_wb_ip7_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7_q_head_r_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_3_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_4_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_5_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_6_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_7_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_8_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_9_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_10_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_11_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_12_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_13_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_14_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_15_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_16_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_17_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_18_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_19_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_20_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_21_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_22_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_23_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_24_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_25_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_26_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_27_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_28_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_29_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_30_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_31_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_32_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_33_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_34_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_35_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_36_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_37_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_38_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_39_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_40_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_41_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_42_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_43_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_44_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_45_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_46_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_47_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_48_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_49_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_50_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_51_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_52_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_53_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_54_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_55_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_56_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_57_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_58_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_59_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_60_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_61_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_62_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_63_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_64_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_65_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_66_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_67_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_68_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_70_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_71_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_72_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_73_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_74_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_75_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_76_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_77_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_78_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_79_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_80_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_81_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_82_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_83_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_84_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_85_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_86_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_87_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_88_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_89_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_90_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_91_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_92_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_93_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_94_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_95_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_96_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_97_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_98_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_99_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_100_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_101_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_102_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_103_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_104_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_105_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_106_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_107_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_108_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_109_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_110_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_111_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_112_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_113_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_114_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_115_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_116_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_117_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_118_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_119_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_120_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_121_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_122_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_123_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_124_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_125_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_126_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_127_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_128_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_129_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_130_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_131_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_132_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7__T_133_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_ip7_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_ip7_q_head_w_en; // @[utils.scala 30:18]
  reg  queue_bits_wb_is_ds [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_15;
  wire  queue_bits_wb_is_ds_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds_q_head_r_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_3_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_4_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_5_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_6_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_7_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_8_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_9_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_10_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_11_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_12_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_13_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_14_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_15_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_16_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_17_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_18_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_19_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_20_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_21_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_22_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_23_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_24_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_25_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_26_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_27_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_28_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_29_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_30_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_31_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_32_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_33_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_34_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_35_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_36_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_37_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_38_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_39_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_40_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_41_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_42_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_43_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_44_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_45_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_46_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_47_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_48_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_49_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_50_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_51_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_52_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_53_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_54_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_55_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_56_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_57_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_58_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_59_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_60_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_61_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_62_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_63_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_64_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_65_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_66_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_67_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_68_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_70_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_71_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_72_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_73_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_74_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_75_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_76_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_77_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_78_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_79_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_80_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_81_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_82_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_83_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_84_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_85_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_86_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_87_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_88_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_89_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_90_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_91_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_92_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_93_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_94_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_95_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_96_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_97_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_98_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_99_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_100_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_101_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_102_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_103_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_104_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_105_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_106_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_107_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_108_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_109_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_110_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_111_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_112_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_113_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_114_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_115_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_116_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_117_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_118_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_119_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_120_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_121_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_122_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_123_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_124_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_125_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_126_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_127_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_128_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_129_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_130_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_131_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_132_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds__T_133_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_ds_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_ds_q_head_w_en; // @[utils.scala 30:18]
  reg  queue_bits_wb_is_br [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_16;
  wire  queue_bits_wb_is_br_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br_q_head_r_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_3_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_4_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_5_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_6_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_7_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_8_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_9_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_10_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_11_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_12_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_13_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_14_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_15_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_16_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_17_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_18_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_19_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_20_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_21_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_22_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_23_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_24_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_25_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_26_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_27_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_28_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_29_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_30_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_31_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_32_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_33_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_34_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_35_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_36_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_37_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_38_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_39_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_40_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_41_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_42_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_43_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_44_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_45_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_46_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_47_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_48_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_49_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_50_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_51_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_52_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_53_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_54_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_55_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_56_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_57_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_58_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_59_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_60_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_61_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_62_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_63_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_64_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_65_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_66_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_67_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_68_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_70_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_71_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_72_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_73_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_74_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_75_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_76_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_77_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_78_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_79_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_80_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_81_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_82_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_83_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_84_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_85_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_86_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_87_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_88_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_89_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_90_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_91_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_92_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_93_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_94_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_95_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_96_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_97_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_98_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_99_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_100_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_101_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_102_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_103_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_104_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_105_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_106_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_107_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_108_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_109_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_110_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_111_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_112_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_113_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_114_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_115_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_116_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_117_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_118_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_119_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_120_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_121_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_122_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_123_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_124_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_125_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_126_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_127_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_128_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_129_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_130_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_131_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_132_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br__T_133_en; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_is_br_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_is_br_q_head_w_en; // @[utils.scala 30:18]
  reg [31:0] queue_bits_wb_npc [0:63]; // @[utils.scala 30:18]
  reg [31:0] _RAND_17;
  wire [31:0] queue_bits_wb_npc_q_head_r_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc_q_head_r_addr; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_3_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_3_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_3_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_3_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_4_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_4_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_4_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_4_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_5_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_5_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_5_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_5_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_6_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_6_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_6_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_6_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_7_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_7_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_7_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_7_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_8_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_8_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_8_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_8_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_9_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_9_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_9_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_9_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_10_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_10_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_10_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_10_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_11_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_11_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_11_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_11_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_12_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_12_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_12_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_12_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_13_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_13_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_13_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_13_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_14_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_14_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_14_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_14_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_15_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_15_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_15_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_15_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_16_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_16_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_16_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_16_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_17_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_17_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_17_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_17_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_18_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_18_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_18_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_18_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_19_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_19_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_19_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_19_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_20_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_20_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_20_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_20_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_21_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_21_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_21_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_21_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_22_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_22_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_22_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_22_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_23_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_23_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_23_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_23_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_24_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_24_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_24_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_24_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_25_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_25_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_25_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_25_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_26_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_26_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_26_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_26_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_27_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_27_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_27_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_27_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_28_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_28_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_28_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_28_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_29_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_29_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_29_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_29_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_30_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_30_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_30_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_30_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_31_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_31_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_31_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_31_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_32_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_32_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_32_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_32_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_33_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_33_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_33_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_33_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_34_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_34_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_34_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_34_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_35_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_35_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_35_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_35_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_36_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_36_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_36_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_36_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_37_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_37_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_37_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_37_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_38_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_38_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_38_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_38_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_39_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_39_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_39_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_39_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_40_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_40_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_40_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_40_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_41_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_41_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_41_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_41_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_42_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_42_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_42_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_42_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_43_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_43_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_43_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_43_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_44_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_44_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_44_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_44_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_45_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_45_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_45_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_45_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_46_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_46_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_46_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_46_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_47_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_47_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_47_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_47_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_48_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_48_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_48_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_48_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_49_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_49_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_49_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_49_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_50_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_50_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_50_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_50_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_51_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_51_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_51_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_51_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_52_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_52_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_52_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_52_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_53_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_53_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_53_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_53_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_54_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_54_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_54_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_54_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_55_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_55_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_55_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_55_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_56_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_56_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_56_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_56_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_57_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_57_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_57_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_57_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_58_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_58_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_58_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_58_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_59_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_59_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_59_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_59_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_60_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_60_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_60_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_60_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_61_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_61_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_61_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_61_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_62_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_62_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_62_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_62_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_63_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_63_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_63_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_63_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_64_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_64_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_64_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_64_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_65_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_65_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_65_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_65_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_66_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_66_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_66_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_66_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_67_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_67_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_67_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_67_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_68_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_68_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_68_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_68_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_70_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_70_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_70_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_70_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_71_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_71_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_71_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_71_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_72_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_72_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_72_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_72_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_73_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_73_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_73_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_73_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_74_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_74_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_74_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_74_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_75_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_75_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_75_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_75_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_76_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_76_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_76_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_76_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_77_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_77_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_77_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_77_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_78_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_78_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_78_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_78_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_79_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_79_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_79_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_79_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_80_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_80_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_80_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_80_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_81_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_81_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_81_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_81_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_82_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_82_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_82_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_82_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_83_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_83_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_83_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_83_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_84_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_84_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_84_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_84_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_85_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_85_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_85_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_85_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_86_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_86_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_86_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_86_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_87_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_87_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_87_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_87_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_88_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_88_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_88_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_88_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_89_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_89_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_89_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_89_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_90_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_90_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_90_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_90_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_91_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_91_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_91_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_91_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_92_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_92_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_92_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_92_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_93_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_93_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_93_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_93_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_94_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_94_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_94_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_94_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_95_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_95_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_95_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_95_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_96_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_96_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_96_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_96_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_97_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_97_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_97_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_97_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_98_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_98_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_98_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_98_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_99_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_99_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_99_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_99_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_100_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_100_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_100_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_100_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_101_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_101_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_101_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_101_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_102_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_102_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_102_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_102_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_103_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_103_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_103_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_103_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_104_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_104_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_104_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_104_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_105_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_105_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_105_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_105_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_106_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_106_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_106_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_106_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_107_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_107_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_107_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_107_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_108_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_108_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_108_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_108_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_109_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_109_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_109_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_109_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_110_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_110_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_110_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_110_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_111_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_111_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_111_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_111_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_112_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_112_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_112_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_112_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_113_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_113_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_113_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_113_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_114_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_114_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_114_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_114_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_115_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_115_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_115_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_115_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_116_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_116_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_116_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_116_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_117_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_117_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_117_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_117_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_118_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_118_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_118_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_118_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_119_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_119_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_119_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_119_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_120_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_120_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_120_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_120_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_121_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_121_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_121_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_121_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_122_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_122_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_122_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_122_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_123_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_123_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_123_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_123_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_124_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_124_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_124_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_124_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_125_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_125_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_125_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_125_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_126_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_126_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_126_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_126_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_127_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_127_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_127_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_127_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_128_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_128_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_128_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_128_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_129_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_129_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_129_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_129_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_130_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_130_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_130_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_130_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_131_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_131_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_131_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_131_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_132_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_132_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_132_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_132_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc__T_133_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc__T_133_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_133_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc__T_133_en; // @[utils.scala 30:18]
  wire [31:0] queue_bits_wb_npc_q_head_w_data; // @[utils.scala 30:18]
  wire [5:0] queue_bits_wb_npc_q_head_w_addr; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc_q_head_w_mask; // @[utils.scala 30:18]
  wire  queue_bits_wb_npc_q_head_w_en; // @[utils.scala 30:18]
  reg [5:0] head; // @[utils.scala 31:21]
  reg [31:0] _RAND_18;
  wire [5:0] _T_2 = head + 6'h1; // @[utils.scala 38:18]
  assign queue_valid_q_head_r_addr = head;
  assign queue_valid_q_head_r_data = queue_valid[queue_valid_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_valid__T_3_data = 1'h1;
  assign queue_valid__T_3_addr = io_enq_0_bits_id;
  assign queue_valid__T_3_mask = 1'h1;
  assign queue_valid__T_3_en = io_enq_0_valid;
  assign queue_valid__T_4_data = 1'h1;
  assign queue_valid__T_4_addr = io_enq_1_bits_id;
  assign queue_valid__T_4_mask = 1'h1;
  assign queue_valid__T_4_en = io_enq_1_valid;
  assign queue_valid__T_5_data = 1'h0;
  assign queue_valid__T_5_addr = 6'h0;
  assign queue_valid__T_5_mask = 1'h1;
  assign queue_valid__T_5_en = 1'h0;
  assign queue_valid__T_6_data = 1'h0;
  assign queue_valid__T_6_addr = 6'h1;
  assign queue_valid__T_6_mask = 1'h1;
  assign queue_valid__T_6_en = 1'h0;
  assign queue_valid__T_7_data = 1'h0;
  assign queue_valid__T_7_addr = 6'h2;
  assign queue_valid__T_7_mask = 1'h1;
  assign queue_valid__T_7_en = 1'h0;
  assign queue_valid__T_8_data = 1'h0;
  assign queue_valid__T_8_addr = 6'h3;
  assign queue_valid__T_8_mask = 1'h1;
  assign queue_valid__T_8_en = 1'h0;
  assign queue_valid__T_9_data = 1'h0;
  assign queue_valid__T_9_addr = 6'h4;
  assign queue_valid__T_9_mask = 1'h1;
  assign queue_valid__T_9_en = 1'h0;
  assign queue_valid__T_10_data = 1'h0;
  assign queue_valid__T_10_addr = 6'h5;
  assign queue_valid__T_10_mask = 1'h1;
  assign queue_valid__T_10_en = 1'h0;
  assign queue_valid__T_11_data = 1'h0;
  assign queue_valid__T_11_addr = 6'h6;
  assign queue_valid__T_11_mask = 1'h1;
  assign queue_valid__T_11_en = 1'h0;
  assign queue_valid__T_12_data = 1'h0;
  assign queue_valid__T_12_addr = 6'h7;
  assign queue_valid__T_12_mask = 1'h1;
  assign queue_valid__T_12_en = 1'h0;
  assign queue_valid__T_13_data = 1'h0;
  assign queue_valid__T_13_addr = 6'h8;
  assign queue_valid__T_13_mask = 1'h1;
  assign queue_valid__T_13_en = 1'h0;
  assign queue_valid__T_14_data = 1'h0;
  assign queue_valid__T_14_addr = 6'h9;
  assign queue_valid__T_14_mask = 1'h1;
  assign queue_valid__T_14_en = 1'h0;
  assign queue_valid__T_15_data = 1'h0;
  assign queue_valid__T_15_addr = 6'ha;
  assign queue_valid__T_15_mask = 1'h1;
  assign queue_valid__T_15_en = 1'h0;
  assign queue_valid__T_16_data = 1'h0;
  assign queue_valid__T_16_addr = 6'hb;
  assign queue_valid__T_16_mask = 1'h1;
  assign queue_valid__T_16_en = 1'h0;
  assign queue_valid__T_17_data = 1'h0;
  assign queue_valid__T_17_addr = 6'hc;
  assign queue_valid__T_17_mask = 1'h1;
  assign queue_valid__T_17_en = 1'h0;
  assign queue_valid__T_18_data = 1'h0;
  assign queue_valid__T_18_addr = 6'hd;
  assign queue_valid__T_18_mask = 1'h1;
  assign queue_valid__T_18_en = 1'h0;
  assign queue_valid__T_19_data = 1'h0;
  assign queue_valid__T_19_addr = 6'he;
  assign queue_valid__T_19_mask = 1'h1;
  assign queue_valid__T_19_en = 1'h0;
  assign queue_valid__T_20_data = 1'h0;
  assign queue_valid__T_20_addr = 6'hf;
  assign queue_valid__T_20_mask = 1'h1;
  assign queue_valid__T_20_en = 1'h0;
  assign queue_valid__T_21_data = 1'h0;
  assign queue_valid__T_21_addr = 6'h10;
  assign queue_valid__T_21_mask = 1'h1;
  assign queue_valid__T_21_en = 1'h0;
  assign queue_valid__T_22_data = 1'h0;
  assign queue_valid__T_22_addr = 6'h11;
  assign queue_valid__T_22_mask = 1'h1;
  assign queue_valid__T_22_en = 1'h0;
  assign queue_valid__T_23_data = 1'h0;
  assign queue_valid__T_23_addr = 6'h12;
  assign queue_valid__T_23_mask = 1'h1;
  assign queue_valid__T_23_en = 1'h0;
  assign queue_valid__T_24_data = 1'h0;
  assign queue_valid__T_24_addr = 6'h13;
  assign queue_valid__T_24_mask = 1'h1;
  assign queue_valid__T_24_en = 1'h0;
  assign queue_valid__T_25_data = 1'h0;
  assign queue_valid__T_25_addr = 6'h14;
  assign queue_valid__T_25_mask = 1'h1;
  assign queue_valid__T_25_en = 1'h0;
  assign queue_valid__T_26_data = 1'h0;
  assign queue_valid__T_26_addr = 6'h15;
  assign queue_valid__T_26_mask = 1'h1;
  assign queue_valid__T_26_en = 1'h0;
  assign queue_valid__T_27_data = 1'h0;
  assign queue_valid__T_27_addr = 6'h16;
  assign queue_valid__T_27_mask = 1'h1;
  assign queue_valid__T_27_en = 1'h0;
  assign queue_valid__T_28_data = 1'h0;
  assign queue_valid__T_28_addr = 6'h17;
  assign queue_valid__T_28_mask = 1'h1;
  assign queue_valid__T_28_en = 1'h0;
  assign queue_valid__T_29_data = 1'h0;
  assign queue_valid__T_29_addr = 6'h18;
  assign queue_valid__T_29_mask = 1'h1;
  assign queue_valid__T_29_en = 1'h0;
  assign queue_valid__T_30_data = 1'h0;
  assign queue_valid__T_30_addr = 6'h19;
  assign queue_valid__T_30_mask = 1'h1;
  assign queue_valid__T_30_en = 1'h0;
  assign queue_valid__T_31_data = 1'h0;
  assign queue_valid__T_31_addr = 6'h1a;
  assign queue_valid__T_31_mask = 1'h1;
  assign queue_valid__T_31_en = 1'h0;
  assign queue_valid__T_32_data = 1'h0;
  assign queue_valid__T_32_addr = 6'h1b;
  assign queue_valid__T_32_mask = 1'h1;
  assign queue_valid__T_32_en = 1'h0;
  assign queue_valid__T_33_data = 1'h0;
  assign queue_valid__T_33_addr = 6'h1c;
  assign queue_valid__T_33_mask = 1'h1;
  assign queue_valid__T_33_en = 1'h0;
  assign queue_valid__T_34_data = 1'h0;
  assign queue_valid__T_34_addr = 6'h1d;
  assign queue_valid__T_34_mask = 1'h1;
  assign queue_valid__T_34_en = 1'h0;
  assign queue_valid__T_35_data = 1'h0;
  assign queue_valid__T_35_addr = 6'h1e;
  assign queue_valid__T_35_mask = 1'h1;
  assign queue_valid__T_35_en = 1'h0;
  assign queue_valid__T_36_data = 1'h0;
  assign queue_valid__T_36_addr = 6'h1f;
  assign queue_valid__T_36_mask = 1'h1;
  assign queue_valid__T_36_en = 1'h0;
  assign queue_valid__T_37_data = 1'h0;
  assign queue_valid__T_37_addr = 6'h20;
  assign queue_valid__T_37_mask = 1'h1;
  assign queue_valid__T_37_en = 1'h0;
  assign queue_valid__T_38_data = 1'h0;
  assign queue_valid__T_38_addr = 6'h21;
  assign queue_valid__T_38_mask = 1'h1;
  assign queue_valid__T_38_en = 1'h0;
  assign queue_valid__T_39_data = 1'h0;
  assign queue_valid__T_39_addr = 6'h22;
  assign queue_valid__T_39_mask = 1'h1;
  assign queue_valid__T_39_en = 1'h0;
  assign queue_valid__T_40_data = 1'h0;
  assign queue_valid__T_40_addr = 6'h23;
  assign queue_valid__T_40_mask = 1'h1;
  assign queue_valid__T_40_en = 1'h0;
  assign queue_valid__T_41_data = 1'h0;
  assign queue_valid__T_41_addr = 6'h24;
  assign queue_valid__T_41_mask = 1'h1;
  assign queue_valid__T_41_en = 1'h0;
  assign queue_valid__T_42_data = 1'h0;
  assign queue_valid__T_42_addr = 6'h25;
  assign queue_valid__T_42_mask = 1'h1;
  assign queue_valid__T_42_en = 1'h0;
  assign queue_valid__T_43_data = 1'h0;
  assign queue_valid__T_43_addr = 6'h26;
  assign queue_valid__T_43_mask = 1'h1;
  assign queue_valid__T_43_en = 1'h0;
  assign queue_valid__T_44_data = 1'h0;
  assign queue_valid__T_44_addr = 6'h27;
  assign queue_valid__T_44_mask = 1'h1;
  assign queue_valid__T_44_en = 1'h0;
  assign queue_valid__T_45_data = 1'h0;
  assign queue_valid__T_45_addr = 6'h28;
  assign queue_valid__T_45_mask = 1'h1;
  assign queue_valid__T_45_en = 1'h0;
  assign queue_valid__T_46_data = 1'h0;
  assign queue_valid__T_46_addr = 6'h29;
  assign queue_valid__T_46_mask = 1'h1;
  assign queue_valid__T_46_en = 1'h0;
  assign queue_valid__T_47_data = 1'h0;
  assign queue_valid__T_47_addr = 6'h2a;
  assign queue_valid__T_47_mask = 1'h1;
  assign queue_valid__T_47_en = 1'h0;
  assign queue_valid__T_48_data = 1'h0;
  assign queue_valid__T_48_addr = 6'h2b;
  assign queue_valid__T_48_mask = 1'h1;
  assign queue_valid__T_48_en = 1'h0;
  assign queue_valid__T_49_data = 1'h0;
  assign queue_valid__T_49_addr = 6'h2c;
  assign queue_valid__T_49_mask = 1'h1;
  assign queue_valid__T_49_en = 1'h0;
  assign queue_valid__T_50_data = 1'h0;
  assign queue_valid__T_50_addr = 6'h2d;
  assign queue_valid__T_50_mask = 1'h1;
  assign queue_valid__T_50_en = 1'h0;
  assign queue_valid__T_51_data = 1'h0;
  assign queue_valid__T_51_addr = 6'h2e;
  assign queue_valid__T_51_mask = 1'h1;
  assign queue_valid__T_51_en = 1'h0;
  assign queue_valid__T_52_data = 1'h0;
  assign queue_valid__T_52_addr = 6'h2f;
  assign queue_valid__T_52_mask = 1'h1;
  assign queue_valid__T_52_en = 1'h0;
  assign queue_valid__T_53_data = 1'h0;
  assign queue_valid__T_53_addr = 6'h30;
  assign queue_valid__T_53_mask = 1'h1;
  assign queue_valid__T_53_en = 1'h0;
  assign queue_valid__T_54_data = 1'h0;
  assign queue_valid__T_54_addr = 6'h31;
  assign queue_valid__T_54_mask = 1'h1;
  assign queue_valid__T_54_en = 1'h0;
  assign queue_valid__T_55_data = 1'h0;
  assign queue_valid__T_55_addr = 6'h32;
  assign queue_valid__T_55_mask = 1'h1;
  assign queue_valid__T_55_en = 1'h0;
  assign queue_valid__T_56_data = 1'h0;
  assign queue_valid__T_56_addr = 6'h33;
  assign queue_valid__T_56_mask = 1'h1;
  assign queue_valid__T_56_en = 1'h0;
  assign queue_valid__T_57_data = 1'h0;
  assign queue_valid__T_57_addr = 6'h34;
  assign queue_valid__T_57_mask = 1'h1;
  assign queue_valid__T_57_en = 1'h0;
  assign queue_valid__T_58_data = 1'h0;
  assign queue_valid__T_58_addr = 6'h35;
  assign queue_valid__T_58_mask = 1'h1;
  assign queue_valid__T_58_en = 1'h0;
  assign queue_valid__T_59_data = 1'h0;
  assign queue_valid__T_59_addr = 6'h36;
  assign queue_valid__T_59_mask = 1'h1;
  assign queue_valid__T_59_en = 1'h0;
  assign queue_valid__T_60_data = 1'h0;
  assign queue_valid__T_60_addr = 6'h37;
  assign queue_valid__T_60_mask = 1'h1;
  assign queue_valid__T_60_en = 1'h0;
  assign queue_valid__T_61_data = 1'h0;
  assign queue_valid__T_61_addr = 6'h38;
  assign queue_valid__T_61_mask = 1'h1;
  assign queue_valid__T_61_en = 1'h0;
  assign queue_valid__T_62_data = 1'h0;
  assign queue_valid__T_62_addr = 6'h39;
  assign queue_valid__T_62_mask = 1'h1;
  assign queue_valid__T_62_en = 1'h0;
  assign queue_valid__T_63_data = 1'h0;
  assign queue_valid__T_63_addr = 6'h3a;
  assign queue_valid__T_63_mask = 1'h1;
  assign queue_valid__T_63_en = 1'h0;
  assign queue_valid__T_64_data = 1'h0;
  assign queue_valid__T_64_addr = 6'h3b;
  assign queue_valid__T_64_mask = 1'h1;
  assign queue_valid__T_64_en = 1'h0;
  assign queue_valid__T_65_data = 1'h0;
  assign queue_valid__T_65_addr = 6'h3c;
  assign queue_valid__T_65_mask = 1'h1;
  assign queue_valid__T_65_en = 1'h0;
  assign queue_valid__T_66_data = 1'h0;
  assign queue_valid__T_66_addr = 6'h3d;
  assign queue_valid__T_66_mask = 1'h1;
  assign queue_valid__T_66_en = 1'h0;
  assign queue_valid__T_67_data = 1'h0;
  assign queue_valid__T_67_addr = 6'h3e;
  assign queue_valid__T_67_mask = 1'h1;
  assign queue_valid__T_67_en = 1'h0;
  assign queue_valid__T_68_data = 1'h0;
  assign queue_valid__T_68_addr = 6'h3f;
  assign queue_valid__T_68_mask = 1'h1;
  assign queue_valid__T_68_en = 1'h0;
  assign queue_valid__T_70_data = 1'h0;
  assign queue_valid__T_70_addr = 6'h0;
  assign queue_valid__T_70_mask = 1'h1;
  assign queue_valid__T_70_en = reset;
  assign queue_valid__T_71_data = 1'h0;
  assign queue_valid__T_71_addr = 6'h1;
  assign queue_valid__T_71_mask = 1'h1;
  assign queue_valid__T_71_en = reset;
  assign queue_valid__T_72_data = 1'h0;
  assign queue_valid__T_72_addr = 6'h2;
  assign queue_valid__T_72_mask = 1'h1;
  assign queue_valid__T_72_en = reset;
  assign queue_valid__T_73_data = 1'h0;
  assign queue_valid__T_73_addr = 6'h3;
  assign queue_valid__T_73_mask = 1'h1;
  assign queue_valid__T_73_en = reset;
  assign queue_valid__T_74_data = 1'h0;
  assign queue_valid__T_74_addr = 6'h4;
  assign queue_valid__T_74_mask = 1'h1;
  assign queue_valid__T_74_en = reset;
  assign queue_valid__T_75_data = 1'h0;
  assign queue_valid__T_75_addr = 6'h5;
  assign queue_valid__T_75_mask = 1'h1;
  assign queue_valid__T_75_en = reset;
  assign queue_valid__T_76_data = 1'h0;
  assign queue_valid__T_76_addr = 6'h6;
  assign queue_valid__T_76_mask = 1'h1;
  assign queue_valid__T_76_en = reset;
  assign queue_valid__T_77_data = 1'h0;
  assign queue_valid__T_77_addr = 6'h7;
  assign queue_valid__T_77_mask = 1'h1;
  assign queue_valid__T_77_en = reset;
  assign queue_valid__T_78_data = 1'h0;
  assign queue_valid__T_78_addr = 6'h8;
  assign queue_valid__T_78_mask = 1'h1;
  assign queue_valid__T_78_en = reset;
  assign queue_valid__T_79_data = 1'h0;
  assign queue_valid__T_79_addr = 6'h9;
  assign queue_valid__T_79_mask = 1'h1;
  assign queue_valid__T_79_en = reset;
  assign queue_valid__T_80_data = 1'h0;
  assign queue_valid__T_80_addr = 6'ha;
  assign queue_valid__T_80_mask = 1'h1;
  assign queue_valid__T_80_en = reset;
  assign queue_valid__T_81_data = 1'h0;
  assign queue_valid__T_81_addr = 6'hb;
  assign queue_valid__T_81_mask = 1'h1;
  assign queue_valid__T_81_en = reset;
  assign queue_valid__T_82_data = 1'h0;
  assign queue_valid__T_82_addr = 6'hc;
  assign queue_valid__T_82_mask = 1'h1;
  assign queue_valid__T_82_en = reset;
  assign queue_valid__T_83_data = 1'h0;
  assign queue_valid__T_83_addr = 6'hd;
  assign queue_valid__T_83_mask = 1'h1;
  assign queue_valid__T_83_en = reset;
  assign queue_valid__T_84_data = 1'h0;
  assign queue_valid__T_84_addr = 6'he;
  assign queue_valid__T_84_mask = 1'h1;
  assign queue_valid__T_84_en = reset;
  assign queue_valid__T_85_data = 1'h0;
  assign queue_valid__T_85_addr = 6'hf;
  assign queue_valid__T_85_mask = 1'h1;
  assign queue_valid__T_85_en = reset;
  assign queue_valid__T_86_data = 1'h0;
  assign queue_valid__T_86_addr = 6'h10;
  assign queue_valid__T_86_mask = 1'h1;
  assign queue_valid__T_86_en = reset;
  assign queue_valid__T_87_data = 1'h0;
  assign queue_valid__T_87_addr = 6'h11;
  assign queue_valid__T_87_mask = 1'h1;
  assign queue_valid__T_87_en = reset;
  assign queue_valid__T_88_data = 1'h0;
  assign queue_valid__T_88_addr = 6'h12;
  assign queue_valid__T_88_mask = 1'h1;
  assign queue_valid__T_88_en = reset;
  assign queue_valid__T_89_data = 1'h0;
  assign queue_valid__T_89_addr = 6'h13;
  assign queue_valid__T_89_mask = 1'h1;
  assign queue_valid__T_89_en = reset;
  assign queue_valid__T_90_data = 1'h0;
  assign queue_valid__T_90_addr = 6'h14;
  assign queue_valid__T_90_mask = 1'h1;
  assign queue_valid__T_90_en = reset;
  assign queue_valid__T_91_data = 1'h0;
  assign queue_valid__T_91_addr = 6'h15;
  assign queue_valid__T_91_mask = 1'h1;
  assign queue_valid__T_91_en = reset;
  assign queue_valid__T_92_data = 1'h0;
  assign queue_valid__T_92_addr = 6'h16;
  assign queue_valid__T_92_mask = 1'h1;
  assign queue_valid__T_92_en = reset;
  assign queue_valid__T_93_data = 1'h0;
  assign queue_valid__T_93_addr = 6'h17;
  assign queue_valid__T_93_mask = 1'h1;
  assign queue_valid__T_93_en = reset;
  assign queue_valid__T_94_data = 1'h0;
  assign queue_valid__T_94_addr = 6'h18;
  assign queue_valid__T_94_mask = 1'h1;
  assign queue_valid__T_94_en = reset;
  assign queue_valid__T_95_data = 1'h0;
  assign queue_valid__T_95_addr = 6'h19;
  assign queue_valid__T_95_mask = 1'h1;
  assign queue_valid__T_95_en = reset;
  assign queue_valid__T_96_data = 1'h0;
  assign queue_valid__T_96_addr = 6'h1a;
  assign queue_valid__T_96_mask = 1'h1;
  assign queue_valid__T_96_en = reset;
  assign queue_valid__T_97_data = 1'h0;
  assign queue_valid__T_97_addr = 6'h1b;
  assign queue_valid__T_97_mask = 1'h1;
  assign queue_valid__T_97_en = reset;
  assign queue_valid__T_98_data = 1'h0;
  assign queue_valid__T_98_addr = 6'h1c;
  assign queue_valid__T_98_mask = 1'h1;
  assign queue_valid__T_98_en = reset;
  assign queue_valid__T_99_data = 1'h0;
  assign queue_valid__T_99_addr = 6'h1d;
  assign queue_valid__T_99_mask = 1'h1;
  assign queue_valid__T_99_en = reset;
  assign queue_valid__T_100_data = 1'h0;
  assign queue_valid__T_100_addr = 6'h1e;
  assign queue_valid__T_100_mask = 1'h1;
  assign queue_valid__T_100_en = reset;
  assign queue_valid__T_101_data = 1'h0;
  assign queue_valid__T_101_addr = 6'h1f;
  assign queue_valid__T_101_mask = 1'h1;
  assign queue_valid__T_101_en = reset;
  assign queue_valid__T_102_data = 1'h0;
  assign queue_valid__T_102_addr = 6'h20;
  assign queue_valid__T_102_mask = 1'h1;
  assign queue_valid__T_102_en = reset;
  assign queue_valid__T_103_data = 1'h0;
  assign queue_valid__T_103_addr = 6'h21;
  assign queue_valid__T_103_mask = 1'h1;
  assign queue_valid__T_103_en = reset;
  assign queue_valid__T_104_data = 1'h0;
  assign queue_valid__T_104_addr = 6'h22;
  assign queue_valid__T_104_mask = 1'h1;
  assign queue_valid__T_104_en = reset;
  assign queue_valid__T_105_data = 1'h0;
  assign queue_valid__T_105_addr = 6'h23;
  assign queue_valid__T_105_mask = 1'h1;
  assign queue_valid__T_105_en = reset;
  assign queue_valid__T_106_data = 1'h0;
  assign queue_valid__T_106_addr = 6'h24;
  assign queue_valid__T_106_mask = 1'h1;
  assign queue_valid__T_106_en = reset;
  assign queue_valid__T_107_data = 1'h0;
  assign queue_valid__T_107_addr = 6'h25;
  assign queue_valid__T_107_mask = 1'h1;
  assign queue_valid__T_107_en = reset;
  assign queue_valid__T_108_data = 1'h0;
  assign queue_valid__T_108_addr = 6'h26;
  assign queue_valid__T_108_mask = 1'h1;
  assign queue_valid__T_108_en = reset;
  assign queue_valid__T_109_data = 1'h0;
  assign queue_valid__T_109_addr = 6'h27;
  assign queue_valid__T_109_mask = 1'h1;
  assign queue_valid__T_109_en = reset;
  assign queue_valid__T_110_data = 1'h0;
  assign queue_valid__T_110_addr = 6'h28;
  assign queue_valid__T_110_mask = 1'h1;
  assign queue_valid__T_110_en = reset;
  assign queue_valid__T_111_data = 1'h0;
  assign queue_valid__T_111_addr = 6'h29;
  assign queue_valid__T_111_mask = 1'h1;
  assign queue_valid__T_111_en = reset;
  assign queue_valid__T_112_data = 1'h0;
  assign queue_valid__T_112_addr = 6'h2a;
  assign queue_valid__T_112_mask = 1'h1;
  assign queue_valid__T_112_en = reset;
  assign queue_valid__T_113_data = 1'h0;
  assign queue_valid__T_113_addr = 6'h2b;
  assign queue_valid__T_113_mask = 1'h1;
  assign queue_valid__T_113_en = reset;
  assign queue_valid__T_114_data = 1'h0;
  assign queue_valid__T_114_addr = 6'h2c;
  assign queue_valid__T_114_mask = 1'h1;
  assign queue_valid__T_114_en = reset;
  assign queue_valid__T_115_data = 1'h0;
  assign queue_valid__T_115_addr = 6'h2d;
  assign queue_valid__T_115_mask = 1'h1;
  assign queue_valid__T_115_en = reset;
  assign queue_valid__T_116_data = 1'h0;
  assign queue_valid__T_116_addr = 6'h2e;
  assign queue_valid__T_116_mask = 1'h1;
  assign queue_valid__T_116_en = reset;
  assign queue_valid__T_117_data = 1'h0;
  assign queue_valid__T_117_addr = 6'h2f;
  assign queue_valid__T_117_mask = 1'h1;
  assign queue_valid__T_117_en = reset;
  assign queue_valid__T_118_data = 1'h0;
  assign queue_valid__T_118_addr = 6'h30;
  assign queue_valid__T_118_mask = 1'h1;
  assign queue_valid__T_118_en = reset;
  assign queue_valid__T_119_data = 1'h0;
  assign queue_valid__T_119_addr = 6'h31;
  assign queue_valid__T_119_mask = 1'h1;
  assign queue_valid__T_119_en = reset;
  assign queue_valid__T_120_data = 1'h0;
  assign queue_valid__T_120_addr = 6'h32;
  assign queue_valid__T_120_mask = 1'h1;
  assign queue_valid__T_120_en = reset;
  assign queue_valid__T_121_data = 1'h0;
  assign queue_valid__T_121_addr = 6'h33;
  assign queue_valid__T_121_mask = 1'h1;
  assign queue_valid__T_121_en = reset;
  assign queue_valid__T_122_data = 1'h0;
  assign queue_valid__T_122_addr = 6'h34;
  assign queue_valid__T_122_mask = 1'h1;
  assign queue_valid__T_122_en = reset;
  assign queue_valid__T_123_data = 1'h0;
  assign queue_valid__T_123_addr = 6'h35;
  assign queue_valid__T_123_mask = 1'h1;
  assign queue_valid__T_123_en = reset;
  assign queue_valid__T_124_data = 1'h0;
  assign queue_valid__T_124_addr = 6'h36;
  assign queue_valid__T_124_mask = 1'h1;
  assign queue_valid__T_124_en = reset;
  assign queue_valid__T_125_data = 1'h0;
  assign queue_valid__T_125_addr = 6'h37;
  assign queue_valid__T_125_mask = 1'h1;
  assign queue_valid__T_125_en = reset;
  assign queue_valid__T_126_data = 1'h0;
  assign queue_valid__T_126_addr = 6'h38;
  assign queue_valid__T_126_mask = 1'h1;
  assign queue_valid__T_126_en = reset;
  assign queue_valid__T_127_data = 1'h0;
  assign queue_valid__T_127_addr = 6'h39;
  assign queue_valid__T_127_mask = 1'h1;
  assign queue_valid__T_127_en = reset;
  assign queue_valid__T_128_data = 1'h0;
  assign queue_valid__T_128_addr = 6'h3a;
  assign queue_valid__T_128_mask = 1'h1;
  assign queue_valid__T_128_en = reset;
  assign queue_valid__T_129_data = 1'h0;
  assign queue_valid__T_129_addr = 6'h3b;
  assign queue_valid__T_129_mask = 1'h1;
  assign queue_valid__T_129_en = reset;
  assign queue_valid__T_130_data = 1'h0;
  assign queue_valid__T_130_addr = 6'h3c;
  assign queue_valid__T_130_mask = 1'h1;
  assign queue_valid__T_130_en = reset;
  assign queue_valid__T_131_data = 1'h0;
  assign queue_valid__T_131_addr = 6'h3d;
  assign queue_valid__T_131_mask = 1'h1;
  assign queue_valid__T_131_en = reset;
  assign queue_valid__T_132_data = 1'h0;
  assign queue_valid__T_132_addr = 6'h3e;
  assign queue_valid__T_132_mask = 1'h1;
  assign queue_valid__T_132_en = reset;
  assign queue_valid__T_133_data = 1'h0;
  assign queue_valid__T_133_addr = 6'h3f;
  assign queue_valid__T_133_mask = 1'h1;
  assign queue_valid__T_133_en = reset;
  assign queue_valid_q_head_w_data = 1'h0;
  assign queue_valid_q_head_w_addr = head;
  assign queue_valid_q_head_w_mask = io_deq_valid;
  assign queue_valid_q_head_w_en = io_deq_valid;
  assign queue_bits_hi_q_head_r_addr = head;
  assign queue_bits_hi_q_head_r_data = queue_bits_hi[queue_bits_hi_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_hi__T_3_data = io_enq_0_bits_data_hi;
  assign queue_bits_hi__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_hi__T_3_mask = 1'h1;
  assign queue_bits_hi__T_3_en = io_enq_0_valid;
  assign queue_bits_hi__T_4_data = io_enq_1_bits_data_hi;
  assign queue_bits_hi__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_hi__T_4_mask = 1'h1;
  assign queue_bits_hi__T_4_en = io_enq_1_valid;
  assign queue_bits_hi__T_5_data = 32'h0;
  assign queue_bits_hi__T_5_addr = 6'h0;
  assign queue_bits_hi__T_5_mask = 1'h0;
  assign queue_bits_hi__T_5_en = 1'h0;
  assign queue_bits_hi__T_6_data = 32'h0;
  assign queue_bits_hi__T_6_addr = 6'h1;
  assign queue_bits_hi__T_6_mask = 1'h0;
  assign queue_bits_hi__T_6_en = 1'h0;
  assign queue_bits_hi__T_7_data = 32'h0;
  assign queue_bits_hi__T_7_addr = 6'h2;
  assign queue_bits_hi__T_7_mask = 1'h0;
  assign queue_bits_hi__T_7_en = 1'h0;
  assign queue_bits_hi__T_8_data = 32'h0;
  assign queue_bits_hi__T_8_addr = 6'h3;
  assign queue_bits_hi__T_8_mask = 1'h0;
  assign queue_bits_hi__T_8_en = 1'h0;
  assign queue_bits_hi__T_9_data = 32'h0;
  assign queue_bits_hi__T_9_addr = 6'h4;
  assign queue_bits_hi__T_9_mask = 1'h0;
  assign queue_bits_hi__T_9_en = 1'h0;
  assign queue_bits_hi__T_10_data = 32'h0;
  assign queue_bits_hi__T_10_addr = 6'h5;
  assign queue_bits_hi__T_10_mask = 1'h0;
  assign queue_bits_hi__T_10_en = 1'h0;
  assign queue_bits_hi__T_11_data = 32'h0;
  assign queue_bits_hi__T_11_addr = 6'h6;
  assign queue_bits_hi__T_11_mask = 1'h0;
  assign queue_bits_hi__T_11_en = 1'h0;
  assign queue_bits_hi__T_12_data = 32'h0;
  assign queue_bits_hi__T_12_addr = 6'h7;
  assign queue_bits_hi__T_12_mask = 1'h0;
  assign queue_bits_hi__T_12_en = 1'h0;
  assign queue_bits_hi__T_13_data = 32'h0;
  assign queue_bits_hi__T_13_addr = 6'h8;
  assign queue_bits_hi__T_13_mask = 1'h0;
  assign queue_bits_hi__T_13_en = 1'h0;
  assign queue_bits_hi__T_14_data = 32'h0;
  assign queue_bits_hi__T_14_addr = 6'h9;
  assign queue_bits_hi__T_14_mask = 1'h0;
  assign queue_bits_hi__T_14_en = 1'h0;
  assign queue_bits_hi__T_15_data = 32'h0;
  assign queue_bits_hi__T_15_addr = 6'ha;
  assign queue_bits_hi__T_15_mask = 1'h0;
  assign queue_bits_hi__T_15_en = 1'h0;
  assign queue_bits_hi__T_16_data = 32'h0;
  assign queue_bits_hi__T_16_addr = 6'hb;
  assign queue_bits_hi__T_16_mask = 1'h0;
  assign queue_bits_hi__T_16_en = 1'h0;
  assign queue_bits_hi__T_17_data = 32'h0;
  assign queue_bits_hi__T_17_addr = 6'hc;
  assign queue_bits_hi__T_17_mask = 1'h0;
  assign queue_bits_hi__T_17_en = 1'h0;
  assign queue_bits_hi__T_18_data = 32'h0;
  assign queue_bits_hi__T_18_addr = 6'hd;
  assign queue_bits_hi__T_18_mask = 1'h0;
  assign queue_bits_hi__T_18_en = 1'h0;
  assign queue_bits_hi__T_19_data = 32'h0;
  assign queue_bits_hi__T_19_addr = 6'he;
  assign queue_bits_hi__T_19_mask = 1'h0;
  assign queue_bits_hi__T_19_en = 1'h0;
  assign queue_bits_hi__T_20_data = 32'h0;
  assign queue_bits_hi__T_20_addr = 6'hf;
  assign queue_bits_hi__T_20_mask = 1'h0;
  assign queue_bits_hi__T_20_en = 1'h0;
  assign queue_bits_hi__T_21_data = 32'h0;
  assign queue_bits_hi__T_21_addr = 6'h10;
  assign queue_bits_hi__T_21_mask = 1'h0;
  assign queue_bits_hi__T_21_en = 1'h0;
  assign queue_bits_hi__T_22_data = 32'h0;
  assign queue_bits_hi__T_22_addr = 6'h11;
  assign queue_bits_hi__T_22_mask = 1'h0;
  assign queue_bits_hi__T_22_en = 1'h0;
  assign queue_bits_hi__T_23_data = 32'h0;
  assign queue_bits_hi__T_23_addr = 6'h12;
  assign queue_bits_hi__T_23_mask = 1'h0;
  assign queue_bits_hi__T_23_en = 1'h0;
  assign queue_bits_hi__T_24_data = 32'h0;
  assign queue_bits_hi__T_24_addr = 6'h13;
  assign queue_bits_hi__T_24_mask = 1'h0;
  assign queue_bits_hi__T_24_en = 1'h0;
  assign queue_bits_hi__T_25_data = 32'h0;
  assign queue_bits_hi__T_25_addr = 6'h14;
  assign queue_bits_hi__T_25_mask = 1'h0;
  assign queue_bits_hi__T_25_en = 1'h0;
  assign queue_bits_hi__T_26_data = 32'h0;
  assign queue_bits_hi__T_26_addr = 6'h15;
  assign queue_bits_hi__T_26_mask = 1'h0;
  assign queue_bits_hi__T_26_en = 1'h0;
  assign queue_bits_hi__T_27_data = 32'h0;
  assign queue_bits_hi__T_27_addr = 6'h16;
  assign queue_bits_hi__T_27_mask = 1'h0;
  assign queue_bits_hi__T_27_en = 1'h0;
  assign queue_bits_hi__T_28_data = 32'h0;
  assign queue_bits_hi__T_28_addr = 6'h17;
  assign queue_bits_hi__T_28_mask = 1'h0;
  assign queue_bits_hi__T_28_en = 1'h0;
  assign queue_bits_hi__T_29_data = 32'h0;
  assign queue_bits_hi__T_29_addr = 6'h18;
  assign queue_bits_hi__T_29_mask = 1'h0;
  assign queue_bits_hi__T_29_en = 1'h0;
  assign queue_bits_hi__T_30_data = 32'h0;
  assign queue_bits_hi__T_30_addr = 6'h19;
  assign queue_bits_hi__T_30_mask = 1'h0;
  assign queue_bits_hi__T_30_en = 1'h0;
  assign queue_bits_hi__T_31_data = 32'h0;
  assign queue_bits_hi__T_31_addr = 6'h1a;
  assign queue_bits_hi__T_31_mask = 1'h0;
  assign queue_bits_hi__T_31_en = 1'h0;
  assign queue_bits_hi__T_32_data = 32'h0;
  assign queue_bits_hi__T_32_addr = 6'h1b;
  assign queue_bits_hi__T_32_mask = 1'h0;
  assign queue_bits_hi__T_32_en = 1'h0;
  assign queue_bits_hi__T_33_data = 32'h0;
  assign queue_bits_hi__T_33_addr = 6'h1c;
  assign queue_bits_hi__T_33_mask = 1'h0;
  assign queue_bits_hi__T_33_en = 1'h0;
  assign queue_bits_hi__T_34_data = 32'h0;
  assign queue_bits_hi__T_34_addr = 6'h1d;
  assign queue_bits_hi__T_34_mask = 1'h0;
  assign queue_bits_hi__T_34_en = 1'h0;
  assign queue_bits_hi__T_35_data = 32'h0;
  assign queue_bits_hi__T_35_addr = 6'h1e;
  assign queue_bits_hi__T_35_mask = 1'h0;
  assign queue_bits_hi__T_35_en = 1'h0;
  assign queue_bits_hi__T_36_data = 32'h0;
  assign queue_bits_hi__T_36_addr = 6'h1f;
  assign queue_bits_hi__T_36_mask = 1'h0;
  assign queue_bits_hi__T_36_en = 1'h0;
  assign queue_bits_hi__T_37_data = 32'h0;
  assign queue_bits_hi__T_37_addr = 6'h20;
  assign queue_bits_hi__T_37_mask = 1'h0;
  assign queue_bits_hi__T_37_en = 1'h0;
  assign queue_bits_hi__T_38_data = 32'h0;
  assign queue_bits_hi__T_38_addr = 6'h21;
  assign queue_bits_hi__T_38_mask = 1'h0;
  assign queue_bits_hi__T_38_en = 1'h0;
  assign queue_bits_hi__T_39_data = 32'h0;
  assign queue_bits_hi__T_39_addr = 6'h22;
  assign queue_bits_hi__T_39_mask = 1'h0;
  assign queue_bits_hi__T_39_en = 1'h0;
  assign queue_bits_hi__T_40_data = 32'h0;
  assign queue_bits_hi__T_40_addr = 6'h23;
  assign queue_bits_hi__T_40_mask = 1'h0;
  assign queue_bits_hi__T_40_en = 1'h0;
  assign queue_bits_hi__T_41_data = 32'h0;
  assign queue_bits_hi__T_41_addr = 6'h24;
  assign queue_bits_hi__T_41_mask = 1'h0;
  assign queue_bits_hi__T_41_en = 1'h0;
  assign queue_bits_hi__T_42_data = 32'h0;
  assign queue_bits_hi__T_42_addr = 6'h25;
  assign queue_bits_hi__T_42_mask = 1'h0;
  assign queue_bits_hi__T_42_en = 1'h0;
  assign queue_bits_hi__T_43_data = 32'h0;
  assign queue_bits_hi__T_43_addr = 6'h26;
  assign queue_bits_hi__T_43_mask = 1'h0;
  assign queue_bits_hi__T_43_en = 1'h0;
  assign queue_bits_hi__T_44_data = 32'h0;
  assign queue_bits_hi__T_44_addr = 6'h27;
  assign queue_bits_hi__T_44_mask = 1'h0;
  assign queue_bits_hi__T_44_en = 1'h0;
  assign queue_bits_hi__T_45_data = 32'h0;
  assign queue_bits_hi__T_45_addr = 6'h28;
  assign queue_bits_hi__T_45_mask = 1'h0;
  assign queue_bits_hi__T_45_en = 1'h0;
  assign queue_bits_hi__T_46_data = 32'h0;
  assign queue_bits_hi__T_46_addr = 6'h29;
  assign queue_bits_hi__T_46_mask = 1'h0;
  assign queue_bits_hi__T_46_en = 1'h0;
  assign queue_bits_hi__T_47_data = 32'h0;
  assign queue_bits_hi__T_47_addr = 6'h2a;
  assign queue_bits_hi__T_47_mask = 1'h0;
  assign queue_bits_hi__T_47_en = 1'h0;
  assign queue_bits_hi__T_48_data = 32'h0;
  assign queue_bits_hi__T_48_addr = 6'h2b;
  assign queue_bits_hi__T_48_mask = 1'h0;
  assign queue_bits_hi__T_48_en = 1'h0;
  assign queue_bits_hi__T_49_data = 32'h0;
  assign queue_bits_hi__T_49_addr = 6'h2c;
  assign queue_bits_hi__T_49_mask = 1'h0;
  assign queue_bits_hi__T_49_en = 1'h0;
  assign queue_bits_hi__T_50_data = 32'h0;
  assign queue_bits_hi__T_50_addr = 6'h2d;
  assign queue_bits_hi__T_50_mask = 1'h0;
  assign queue_bits_hi__T_50_en = 1'h0;
  assign queue_bits_hi__T_51_data = 32'h0;
  assign queue_bits_hi__T_51_addr = 6'h2e;
  assign queue_bits_hi__T_51_mask = 1'h0;
  assign queue_bits_hi__T_51_en = 1'h0;
  assign queue_bits_hi__T_52_data = 32'h0;
  assign queue_bits_hi__T_52_addr = 6'h2f;
  assign queue_bits_hi__T_52_mask = 1'h0;
  assign queue_bits_hi__T_52_en = 1'h0;
  assign queue_bits_hi__T_53_data = 32'h0;
  assign queue_bits_hi__T_53_addr = 6'h30;
  assign queue_bits_hi__T_53_mask = 1'h0;
  assign queue_bits_hi__T_53_en = 1'h0;
  assign queue_bits_hi__T_54_data = 32'h0;
  assign queue_bits_hi__T_54_addr = 6'h31;
  assign queue_bits_hi__T_54_mask = 1'h0;
  assign queue_bits_hi__T_54_en = 1'h0;
  assign queue_bits_hi__T_55_data = 32'h0;
  assign queue_bits_hi__T_55_addr = 6'h32;
  assign queue_bits_hi__T_55_mask = 1'h0;
  assign queue_bits_hi__T_55_en = 1'h0;
  assign queue_bits_hi__T_56_data = 32'h0;
  assign queue_bits_hi__T_56_addr = 6'h33;
  assign queue_bits_hi__T_56_mask = 1'h0;
  assign queue_bits_hi__T_56_en = 1'h0;
  assign queue_bits_hi__T_57_data = 32'h0;
  assign queue_bits_hi__T_57_addr = 6'h34;
  assign queue_bits_hi__T_57_mask = 1'h0;
  assign queue_bits_hi__T_57_en = 1'h0;
  assign queue_bits_hi__T_58_data = 32'h0;
  assign queue_bits_hi__T_58_addr = 6'h35;
  assign queue_bits_hi__T_58_mask = 1'h0;
  assign queue_bits_hi__T_58_en = 1'h0;
  assign queue_bits_hi__T_59_data = 32'h0;
  assign queue_bits_hi__T_59_addr = 6'h36;
  assign queue_bits_hi__T_59_mask = 1'h0;
  assign queue_bits_hi__T_59_en = 1'h0;
  assign queue_bits_hi__T_60_data = 32'h0;
  assign queue_bits_hi__T_60_addr = 6'h37;
  assign queue_bits_hi__T_60_mask = 1'h0;
  assign queue_bits_hi__T_60_en = 1'h0;
  assign queue_bits_hi__T_61_data = 32'h0;
  assign queue_bits_hi__T_61_addr = 6'h38;
  assign queue_bits_hi__T_61_mask = 1'h0;
  assign queue_bits_hi__T_61_en = 1'h0;
  assign queue_bits_hi__T_62_data = 32'h0;
  assign queue_bits_hi__T_62_addr = 6'h39;
  assign queue_bits_hi__T_62_mask = 1'h0;
  assign queue_bits_hi__T_62_en = 1'h0;
  assign queue_bits_hi__T_63_data = 32'h0;
  assign queue_bits_hi__T_63_addr = 6'h3a;
  assign queue_bits_hi__T_63_mask = 1'h0;
  assign queue_bits_hi__T_63_en = 1'h0;
  assign queue_bits_hi__T_64_data = 32'h0;
  assign queue_bits_hi__T_64_addr = 6'h3b;
  assign queue_bits_hi__T_64_mask = 1'h0;
  assign queue_bits_hi__T_64_en = 1'h0;
  assign queue_bits_hi__T_65_data = 32'h0;
  assign queue_bits_hi__T_65_addr = 6'h3c;
  assign queue_bits_hi__T_65_mask = 1'h0;
  assign queue_bits_hi__T_65_en = 1'h0;
  assign queue_bits_hi__T_66_data = 32'h0;
  assign queue_bits_hi__T_66_addr = 6'h3d;
  assign queue_bits_hi__T_66_mask = 1'h0;
  assign queue_bits_hi__T_66_en = 1'h0;
  assign queue_bits_hi__T_67_data = 32'h0;
  assign queue_bits_hi__T_67_addr = 6'h3e;
  assign queue_bits_hi__T_67_mask = 1'h0;
  assign queue_bits_hi__T_67_en = 1'h0;
  assign queue_bits_hi__T_68_data = 32'h0;
  assign queue_bits_hi__T_68_addr = 6'h3f;
  assign queue_bits_hi__T_68_mask = 1'h0;
  assign queue_bits_hi__T_68_en = 1'h0;
  assign queue_bits_hi__T_70_data = 32'h0;
  assign queue_bits_hi__T_70_addr = 6'h0;
  assign queue_bits_hi__T_70_mask = 1'h0;
  assign queue_bits_hi__T_70_en = reset;
  assign queue_bits_hi__T_71_data = 32'h0;
  assign queue_bits_hi__T_71_addr = 6'h1;
  assign queue_bits_hi__T_71_mask = 1'h0;
  assign queue_bits_hi__T_71_en = reset;
  assign queue_bits_hi__T_72_data = 32'h0;
  assign queue_bits_hi__T_72_addr = 6'h2;
  assign queue_bits_hi__T_72_mask = 1'h0;
  assign queue_bits_hi__T_72_en = reset;
  assign queue_bits_hi__T_73_data = 32'h0;
  assign queue_bits_hi__T_73_addr = 6'h3;
  assign queue_bits_hi__T_73_mask = 1'h0;
  assign queue_bits_hi__T_73_en = reset;
  assign queue_bits_hi__T_74_data = 32'h0;
  assign queue_bits_hi__T_74_addr = 6'h4;
  assign queue_bits_hi__T_74_mask = 1'h0;
  assign queue_bits_hi__T_74_en = reset;
  assign queue_bits_hi__T_75_data = 32'h0;
  assign queue_bits_hi__T_75_addr = 6'h5;
  assign queue_bits_hi__T_75_mask = 1'h0;
  assign queue_bits_hi__T_75_en = reset;
  assign queue_bits_hi__T_76_data = 32'h0;
  assign queue_bits_hi__T_76_addr = 6'h6;
  assign queue_bits_hi__T_76_mask = 1'h0;
  assign queue_bits_hi__T_76_en = reset;
  assign queue_bits_hi__T_77_data = 32'h0;
  assign queue_bits_hi__T_77_addr = 6'h7;
  assign queue_bits_hi__T_77_mask = 1'h0;
  assign queue_bits_hi__T_77_en = reset;
  assign queue_bits_hi__T_78_data = 32'h0;
  assign queue_bits_hi__T_78_addr = 6'h8;
  assign queue_bits_hi__T_78_mask = 1'h0;
  assign queue_bits_hi__T_78_en = reset;
  assign queue_bits_hi__T_79_data = 32'h0;
  assign queue_bits_hi__T_79_addr = 6'h9;
  assign queue_bits_hi__T_79_mask = 1'h0;
  assign queue_bits_hi__T_79_en = reset;
  assign queue_bits_hi__T_80_data = 32'h0;
  assign queue_bits_hi__T_80_addr = 6'ha;
  assign queue_bits_hi__T_80_mask = 1'h0;
  assign queue_bits_hi__T_80_en = reset;
  assign queue_bits_hi__T_81_data = 32'h0;
  assign queue_bits_hi__T_81_addr = 6'hb;
  assign queue_bits_hi__T_81_mask = 1'h0;
  assign queue_bits_hi__T_81_en = reset;
  assign queue_bits_hi__T_82_data = 32'h0;
  assign queue_bits_hi__T_82_addr = 6'hc;
  assign queue_bits_hi__T_82_mask = 1'h0;
  assign queue_bits_hi__T_82_en = reset;
  assign queue_bits_hi__T_83_data = 32'h0;
  assign queue_bits_hi__T_83_addr = 6'hd;
  assign queue_bits_hi__T_83_mask = 1'h0;
  assign queue_bits_hi__T_83_en = reset;
  assign queue_bits_hi__T_84_data = 32'h0;
  assign queue_bits_hi__T_84_addr = 6'he;
  assign queue_bits_hi__T_84_mask = 1'h0;
  assign queue_bits_hi__T_84_en = reset;
  assign queue_bits_hi__T_85_data = 32'h0;
  assign queue_bits_hi__T_85_addr = 6'hf;
  assign queue_bits_hi__T_85_mask = 1'h0;
  assign queue_bits_hi__T_85_en = reset;
  assign queue_bits_hi__T_86_data = 32'h0;
  assign queue_bits_hi__T_86_addr = 6'h10;
  assign queue_bits_hi__T_86_mask = 1'h0;
  assign queue_bits_hi__T_86_en = reset;
  assign queue_bits_hi__T_87_data = 32'h0;
  assign queue_bits_hi__T_87_addr = 6'h11;
  assign queue_bits_hi__T_87_mask = 1'h0;
  assign queue_bits_hi__T_87_en = reset;
  assign queue_bits_hi__T_88_data = 32'h0;
  assign queue_bits_hi__T_88_addr = 6'h12;
  assign queue_bits_hi__T_88_mask = 1'h0;
  assign queue_bits_hi__T_88_en = reset;
  assign queue_bits_hi__T_89_data = 32'h0;
  assign queue_bits_hi__T_89_addr = 6'h13;
  assign queue_bits_hi__T_89_mask = 1'h0;
  assign queue_bits_hi__T_89_en = reset;
  assign queue_bits_hi__T_90_data = 32'h0;
  assign queue_bits_hi__T_90_addr = 6'h14;
  assign queue_bits_hi__T_90_mask = 1'h0;
  assign queue_bits_hi__T_90_en = reset;
  assign queue_bits_hi__T_91_data = 32'h0;
  assign queue_bits_hi__T_91_addr = 6'h15;
  assign queue_bits_hi__T_91_mask = 1'h0;
  assign queue_bits_hi__T_91_en = reset;
  assign queue_bits_hi__T_92_data = 32'h0;
  assign queue_bits_hi__T_92_addr = 6'h16;
  assign queue_bits_hi__T_92_mask = 1'h0;
  assign queue_bits_hi__T_92_en = reset;
  assign queue_bits_hi__T_93_data = 32'h0;
  assign queue_bits_hi__T_93_addr = 6'h17;
  assign queue_bits_hi__T_93_mask = 1'h0;
  assign queue_bits_hi__T_93_en = reset;
  assign queue_bits_hi__T_94_data = 32'h0;
  assign queue_bits_hi__T_94_addr = 6'h18;
  assign queue_bits_hi__T_94_mask = 1'h0;
  assign queue_bits_hi__T_94_en = reset;
  assign queue_bits_hi__T_95_data = 32'h0;
  assign queue_bits_hi__T_95_addr = 6'h19;
  assign queue_bits_hi__T_95_mask = 1'h0;
  assign queue_bits_hi__T_95_en = reset;
  assign queue_bits_hi__T_96_data = 32'h0;
  assign queue_bits_hi__T_96_addr = 6'h1a;
  assign queue_bits_hi__T_96_mask = 1'h0;
  assign queue_bits_hi__T_96_en = reset;
  assign queue_bits_hi__T_97_data = 32'h0;
  assign queue_bits_hi__T_97_addr = 6'h1b;
  assign queue_bits_hi__T_97_mask = 1'h0;
  assign queue_bits_hi__T_97_en = reset;
  assign queue_bits_hi__T_98_data = 32'h0;
  assign queue_bits_hi__T_98_addr = 6'h1c;
  assign queue_bits_hi__T_98_mask = 1'h0;
  assign queue_bits_hi__T_98_en = reset;
  assign queue_bits_hi__T_99_data = 32'h0;
  assign queue_bits_hi__T_99_addr = 6'h1d;
  assign queue_bits_hi__T_99_mask = 1'h0;
  assign queue_bits_hi__T_99_en = reset;
  assign queue_bits_hi__T_100_data = 32'h0;
  assign queue_bits_hi__T_100_addr = 6'h1e;
  assign queue_bits_hi__T_100_mask = 1'h0;
  assign queue_bits_hi__T_100_en = reset;
  assign queue_bits_hi__T_101_data = 32'h0;
  assign queue_bits_hi__T_101_addr = 6'h1f;
  assign queue_bits_hi__T_101_mask = 1'h0;
  assign queue_bits_hi__T_101_en = reset;
  assign queue_bits_hi__T_102_data = 32'h0;
  assign queue_bits_hi__T_102_addr = 6'h20;
  assign queue_bits_hi__T_102_mask = 1'h0;
  assign queue_bits_hi__T_102_en = reset;
  assign queue_bits_hi__T_103_data = 32'h0;
  assign queue_bits_hi__T_103_addr = 6'h21;
  assign queue_bits_hi__T_103_mask = 1'h0;
  assign queue_bits_hi__T_103_en = reset;
  assign queue_bits_hi__T_104_data = 32'h0;
  assign queue_bits_hi__T_104_addr = 6'h22;
  assign queue_bits_hi__T_104_mask = 1'h0;
  assign queue_bits_hi__T_104_en = reset;
  assign queue_bits_hi__T_105_data = 32'h0;
  assign queue_bits_hi__T_105_addr = 6'h23;
  assign queue_bits_hi__T_105_mask = 1'h0;
  assign queue_bits_hi__T_105_en = reset;
  assign queue_bits_hi__T_106_data = 32'h0;
  assign queue_bits_hi__T_106_addr = 6'h24;
  assign queue_bits_hi__T_106_mask = 1'h0;
  assign queue_bits_hi__T_106_en = reset;
  assign queue_bits_hi__T_107_data = 32'h0;
  assign queue_bits_hi__T_107_addr = 6'h25;
  assign queue_bits_hi__T_107_mask = 1'h0;
  assign queue_bits_hi__T_107_en = reset;
  assign queue_bits_hi__T_108_data = 32'h0;
  assign queue_bits_hi__T_108_addr = 6'h26;
  assign queue_bits_hi__T_108_mask = 1'h0;
  assign queue_bits_hi__T_108_en = reset;
  assign queue_bits_hi__T_109_data = 32'h0;
  assign queue_bits_hi__T_109_addr = 6'h27;
  assign queue_bits_hi__T_109_mask = 1'h0;
  assign queue_bits_hi__T_109_en = reset;
  assign queue_bits_hi__T_110_data = 32'h0;
  assign queue_bits_hi__T_110_addr = 6'h28;
  assign queue_bits_hi__T_110_mask = 1'h0;
  assign queue_bits_hi__T_110_en = reset;
  assign queue_bits_hi__T_111_data = 32'h0;
  assign queue_bits_hi__T_111_addr = 6'h29;
  assign queue_bits_hi__T_111_mask = 1'h0;
  assign queue_bits_hi__T_111_en = reset;
  assign queue_bits_hi__T_112_data = 32'h0;
  assign queue_bits_hi__T_112_addr = 6'h2a;
  assign queue_bits_hi__T_112_mask = 1'h0;
  assign queue_bits_hi__T_112_en = reset;
  assign queue_bits_hi__T_113_data = 32'h0;
  assign queue_bits_hi__T_113_addr = 6'h2b;
  assign queue_bits_hi__T_113_mask = 1'h0;
  assign queue_bits_hi__T_113_en = reset;
  assign queue_bits_hi__T_114_data = 32'h0;
  assign queue_bits_hi__T_114_addr = 6'h2c;
  assign queue_bits_hi__T_114_mask = 1'h0;
  assign queue_bits_hi__T_114_en = reset;
  assign queue_bits_hi__T_115_data = 32'h0;
  assign queue_bits_hi__T_115_addr = 6'h2d;
  assign queue_bits_hi__T_115_mask = 1'h0;
  assign queue_bits_hi__T_115_en = reset;
  assign queue_bits_hi__T_116_data = 32'h0;
  assign queue_bits_hi__T_116_addr = 6'h2e;
  assign queue_bits_hi__T_116_mask = 1'h0;
  assign queue_bits_hi__T_116_en = reset;
  assign queue_bits_hi__T_117_data = 32'h0;
  assign queue_bits_hi__T_117_addr = 6'h2f;
  assign queue_bits_hi__T_117_mask = 1'h0;
  assign queue_bits_hi__T_117_en = reset;
  assign queue_bits_hi__T_118_data = 32'h0;
  assign queue_bits_hi__T_118_addr = 6'h30;
  assign queue_bits_hi__T_118_mask = 1'h0;
  assign queue_bits_hi__T_118_en = reset;
  assign queue_bits_hi__T_119_data = 32'h0;
  assign queue_bits_hi__T_119_addr = 6'h31;
  assign queue_bits_hi__T_119_mask = 1'h0;
  assign queue_bits_hi__T_119_en = reset;
  assign queue_bits_hi__T_120_data = 32'h0;
  assign queue_bits_hi__T_120_addr = 6'h32;
  assign queue_bits_hi__T_120_mask = 1'h0;
  assign queue_bits_hi__T_120_en = reset;
  assign queue_bits_hi__T_121_data = 32'h0;
  assign queue_bits_hi__T_121_addr = 6'h33;
  assign queue_bits_hi__T_121_mask = 1'h0;
  assign queue_bits_hi__T_121_en = reset;
  assign queue_bits_hi__T_122_data = 32'h0;
  assign queue_bits_hi__T_122_addr = 6'h34;
  assign queue_bits_hi__T_122_mask = 1'h0;
  assign queue_bits_hi__T_122_en = reset;
  assign queue_bits_hi__T_123_data = 32'h0;
  assign queue_bits_hi__T_123_addr = 6'h35;
  assign queue_bits_hi__T_123_mask = 1'h0;
  assign queue_bits_hi__T_123_en = reset;
  assign queue_bits_hi__T_124_data = 32'h0;
  assign queue_bits_hi__T_124_addr = 6'h36;
  assign queue_bits_hi__T_124_mask = 1'h0;
  assign queue_bits_hi__T_124_en = reset;
  assign queue_bits_hi__T_125_data = 32'h0;
  assign queue_bits_hi__T_125_addr = 6'h37;
  assign queue_bits_hi__T_125_mask = 1'h0;
  assign queue_bits_hi__T_125_en = reset;
  assign queue_bits_hi__T_126_data = 32'h0;
  assign queue_bits_hi__T_126_addr = 6'h38;
  assign queue_bits_hi__T_126_mask = 1'h0;
  assign queue_bits_hi__T_126_en = reset;
  assign queue_bits_hi__T_127_data = 32'h0;
  assign queue_bits_hi__T_127_addr = 6'h39;
  assign queue_bits_hi__T_127_mask = 1'h0;
  assign queue_bits_hi__T_127_en = reset;
  assign queue_bits_hi__T_128_data = 32'h0;
  assign queue_bits_hi__T_128_addr = 6'h3a;
  assign queue_bits_hi__T_128_mask = 1'h0;
  assign queue_bits_hi__T_128_en = reset;
  assign queue_bits_hi__T_129_data = 32'h0;
  assign queue_bits_hi__T_129_addr = 6'h3b;
  assign queue_bits_hi__T_129_mask = 1'h0;
  assign queue_bits_hi__T_129_en = reset;
  assign queue_bits_hi__T_130_data = 32'h0;
  assign queue_bits_hi__T_130_addr = 6'h3c;
  assign queue_bits_hi__T_130_mask = 1'h0;
  assign queue_bits_hi__T_130_en = reset;
  assign queue_bits_hi__T_131_data = 32'h0;
  assign queue_bits_hi__T_131_addr = 6'h3d;
  assign queue_bits_hi__T_131_mask = 1'h0;
  assign queue_bits_hi__T_131_en = reset;
  assign queue_bits_hi__T_132_data = 32'h0;
  assign queue_bits_hi__T_132_addr = 6'h3e;
  assign queue_bits_hi__T_132_mask = 1'h0;
  assign queue_bits_hi__T_132_en = reset;
  assign queue_bits_hi__T_133_data = 32'h0;
  assign queue_bits_hi__T_133_addr = 6'h3f;
  assign queue_bits_hi__T_133_mask = 1'h0;
  assign queue_bits_hi__T_133_en = reset;
  assign queue_bits_hi_q_head_w_data = 32'h0;
  assign queue_bits_hi_q_head_w_addr = head;
  assign queue_bits_hi_q_head_w_mask = 1'h0;
  assign queue_bits_hi_q_head_w_en = io_deq_valid;
  assign queue_bits_lo_q_head_r_addr = head;
  assign queue_bits_lo_q_head_r_data = queue_bits_lo[queue_bits_lo_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_lo__T_3_data = io_enq_0_bits_data_lo;
  assign queue_bits_lo__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_lo__T_3_mask = 1'h1;
  assign queue_bits_lo__T_3_en = io_enq_0_valid;
  assign queue_bits_lo__T_4_data = io_enq_1_bits_data_lo;
  assign queue_bits_lo__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_lo__T_4_mask = 1'h1;
  assign queue_bits_lo__T_4_en = io_enq_1_valid;
  assign queue_bits_lo__T_5_data = 32'h0;
  assign queue_bits_lo__T_5_addr = 6'h0;
  assign queue_bits_lo__T_5_mask = 1'h0;
  assign queue_bits_lo__T_5_en = 1'h0;
  assign queue_bits_lo__T_6_data = 32'h0;
  assign queue_bits_lo__T_6_addr = 6'h1;
  assign queue_bits_lo__T_6_mask = 1'h0;
  assign queue_bits_lo__T_6_en = 1'h0;
  assign queue_bits_lo__T_7_data = 32'h0;
  assign queue_bits_lo__T_7_addr = 6'h2;
  assign queue_bits_lo__T_7_mask = 1'h0;
  assign queue_bits_lo__T_7_en = 1'h0;
  assign queue_bits_lo__T_8_data = 32'h0;
  assign queue_bits_lo__T_8_addr = 6'h3;
  assign queue_bits_lo__T_8_mask = 1'h0;
  assign queue_bits_lo__T_8_en = 1'h0;
  assign queue_bits_lo__T_9_data = 32'h0;
  assign queue_bits_lo__T_9_addr = 6'h4;
  assign queue_bits_lo__T_9_mask = 1'h0;
  assign queue_bits_lo__T_9_en = 1'h0;
  assign queue_bits_lo__T_10_data = 32'h0;
  assign queue_bits_lo__T_10_addr = 6'h5;
  assign queue_bits_lo__T_10_mask = 1'h0;
  assign queue_bits_lo__T_10_en = 1'h0;
  assign queue_bits_lo__T_11_data = 32'h0;
  assign queue_bits_lo__T_11_addr = 6'h6;
  assign queue_bits_lo__T_11_mask = 1'h0;
  assign queue_bits_lo__T_11_en = 1'h0;
  assign queue_bits_lo__T_12_data = 32'h0;
  assign queue_bits_lo__T_12_addr = 6'h7;
  assign queue_bits_lo__T_12_mask = 1'h0;
  assign queue_bits_lo__T_12_en = 1'h0;
  assign queue_bits_lo__T_13_data = 32'h0;
  assign queue_bits_lo__T_13_addr = 6'h8;
  assign queue_bits_lo__T_13_mask = 1'h0;
  assign queue_bits_lo__T_13_en = 1'h0;
  assign queue_bits_lo__T_14_data = 32'h0;
  assign queue_bits_lo__T_14_addr = 6'h9;
  assign queue_bits_lo__T_14_mask = 1'h0;
  assign queue_bits_lo__T_14_en = 1'h0;
  assign queue_bits_lo__T_15_data = 32'h0;
  assign queue_bits_lo__T_15_addr = 6'ha;
  assign queue_bits_lo__T_15_mask = 1'h0;
  assign queue_bits_lo__T_15_en = 1'h0;
  assign queue_bits_lo__T_16_data = 32'h0;
  assign queue_bits_lo__T_16_addr = 6'hb;
  assign queue_bits_lo__T_16_mask = 1'h0;
  assign queue_bits_lo__T_16_en = 1'h0;
  assign queue_bits_lo__T_17_data = 32'h0;
  assign queue_bits_lo__T_17_addr = 6'hc;
  assign queue_bits_lo__T_17_mask = 1'h0;
  assign queue_bits_lo__T_17_en = 1'h0;
  assign queue_bits_lo__T_18_data = 32'h0;
  assign queue_bits_lo__T_18_addr = 6'hd;
  assign queue_bits_lo__T_18_mask = 1'h0;
  assign queue_bits_lo__T_18_en = 1'h0;
  assign queue_bits_lo__T_19_data = 32'h0;
  assign queue_bits_lo__T_19_addr = 6'he;
  assign queue_bits_lo__T_19_mask = 1'h0;
  assign queue_bits_lo__T_19_en = 1'h0;
  assign queue_bits_lo__T_20_data = 32'h0;
  assign queue_bits_lo__T_20_addr = 6'hf;
  assign queue_bits_lo__T_20_mask = 1'h0;
  assign queue_bits_lo__T_20_en = 1'h0;
  assign queue_bits_lo__T_21_data = 32'h0;
  assign queue_bits_lo__T_21_addr = 6'h10;
  assign queue_bits_lo__T_21_mask = 1'h0;
  assign queue_bits_lo__T_21_en = 1'h0;
  assign queue_bits_lo__T_22_data = 32'h0;
  assign queue_bits_lo__T_22_addr = 6'h11;
  assign queue_bits_lo__T_22_mask = 1'h0;
  assign queue_bits_lo__T_22_en = 1'h0;
  assign queue_bits_lo__T_23_data = 32'h0;
  assign queue_bits_lo__T_23_addr = 6'h12;
  assign queue_bits_lo__T_23_mask = 1'h0;
  assign queue_bits_lo__T_23_en = 1'h0;
  assign queue_bits_lo__T_24_data = 32'h0;
  assign queue_bits_lo__T_24_addr = 6'h13;
  assign queue_bits_lo__T_24_mask = 1'h0;
  assign queue_bits_lo__T_24_en = 1'h0;
  assign queue_bits_lo__T_25_data = 32'h0;
  assign queue_bits_lo__T_25_addr = 6'h14;
  assign queue_bits_lo__T_25_mask = 1'h0;
  assign queue_bits_lo__T_25_en = 1'h0;
  assign queue_bits_lo__T_26_data = 32'h0;
  assign queue_bits_lo__T_26_addr = 6'h15;
  assign queue_bits_lo__T_26_mask = 1'h0;
  assign queue_bits_lo__T_26_en = 1'h0;
  assign queue_bits_lo__T_27_data = 32'h0;
  assign queue_bits_lo__T_27_addr = 6'h16;
  assign queue_bits_lo__T_27_mask = 1'h0;
  assign queue_bits_lo__T_27_en = 1'h0;
  assign queue_bits_lo__T_28_data = 32'h0;
  assign queue_bits_lo__T_28_addr = 6'h17;
  assign queue_bits_lo__T_28_mask = 1'h0;
  assign queue_bits_lo__T_28_en = 1'h0;
  assign queue_bits_lo__T_29_data = 32'h0;
  assign queue_bits_lo__T_29_addr = 6'h18;
  assign queue_bits_lo__T_29_mask = 1'h0;
  assign queue_bits_lo__T_29_en = 1'h0;
  assign queue_bits_lo__T_30_data = 32'h0;
  assign queue_bits_lo__T_30_addr = 6'h19;
  assign queue_bits_lo__T_30_mask = 1'h0;
  assign queue_bits_lo__T_30_en = 1'h0;
  assign queue_bits_lo__T_31_data = 32'h0;
  assign queue_bits_lo__T_31_addr = 6'h1a;
  assign queue_bits_lo__T_31_mask = 1'h0;
  assign queue_bits_lo__T_31_en = 1'h0;
  assign queue_bits_lo__T_32_data = 32'h0;
  assign queue_bits_lo__T_32_addr = 6'h1b;
  assign queue_bits_lo__T_32_mask = 1'h0;
  assign queue_bits_lo__T_32_en = 1'h0;
  assign queue_bits_lo__T_33_data = 32'h0;
  assign queue_bits_lo__T_33_addr = 6'h1c;
  assign queue_bits_lo__T_33_mask = 1'h0;
  assign queue_bits_lo__T_33_en = 1'h0;
  assign queue_bits_lo__T_34_data = 32'h0;
  assign queue_bits_lo__T_34_addr = 6'h1d;
  assign queue_bits_lo__T_34_mask = 1'h0;
  assign queue_bits_lo__T_34_en = 1'h0;
  assign queue_bits_lo__T_35_data = 32'h0;
  assign queue_bits_lo__T_35_addr = 6'h1e;
  assign queue_bits_lo__T_35_mask = 1'h0;
  assign queue_bits_lo__T_35_en = 1'h0;
  assign queue_bits_lo__T_36_data = 32'h0;
  assign queue_bits_lo__T_36_addr = 6'h1f;
  assign queue_bits_lo__T_36_mask = 1'h0;
  assign queue_bits_lo__T_36_en = 1'h0;
  assign queue_bits_lo__T_37_data = 32'h0;
  assign queue_bits_lo__T_37_addr = 6'h20;
  assign queue_bits_lo__T_37_mask = 1'h0;
  assign queue_bits_lo__T_37_en = 1'h0;
  assign queue_bits_lo__T_38_data = 32'h0;
  assign queue_bits_lo__T_38_addr = 6'h21;
  assign queue_bits_lo__T_38_mask = 1'h0;
  assign queue_bits_lo__T_38_en = 1'h0;
  assign queue_bits_lo__T_39_data = 32'h0;
  assign queue_bits_lo__T_39_addr = 6'h22;
  assign queue_bits_lo__T_39_mask = 1'h0;
  assign queue_bits_lo__T_39_en = 1'h0;
  assign queue_bits_lo__T_40_data = 32'h0;
  assign queue_bits_lo__T_40_addr = 6'h23;
  assign queue_bits_lo__T_40_mask = 1'h0;
  assign queue_bits_lo__T_40_en = 1'h0;
  assign queue_bits_lo__T_41_data = 32'h0;
  assign queue_bits_lo__T_41_addr = 6'h24;
  assign queue_bits_lo__T_41_mask = 1'h0;
  assign queue_bits_lo__T_41_en = 1'h0;
  assign queue_bits_lo__T_42_data = 32'h0;
  assign queue_bits_lo__T_42_addr = 6'h25;
  assign queue_bits_lo__T_42_mask = 1'h0;
  assign queue_bits_lo__T_42_en = 1'h0;
  assign queue_bits_lo__T_43_data = 32'h0;
  assign queue_bits_lo__T_43_addr = 6'h26;
  assign queue_bits_lo__T_43_mask = 1'h0;
  assign queue_bits_lo__T_43_en = 1'h0;
  assign queue_bits_lo__T_44_data = 32'h0;
  assign queue_bits_lo__T_44_addr = 6'h27;
  assign queue_bits_lo__T_44_mask = 1'h0;
  assign queue_bits_lo__T_44_en = 1'h0;
  assign queue_bits_lo__T_45_data = 32'h0;
  assign queue_bits_lo__T_45_addr = 6'h28;
  assign queue_bits_lo__T_45_mask = 1'h0;
  assign queue_bits_lo__T_45_en = 1'h0;
  assign queue_bits_lo__T_46_data = 32'h0;
  assign queue_bits_lo__T_46_addr = 6'h29;
  assign queue_bits_lo__T_46_mask = 1'h0;
  assign queue_bits_lo__T_46_en = 1'h0;
  assign queue_bits_lo__T_47_data = 32'h0;
  assign queue_bits_lo__T_47_addr = 6'h2a;
  assign queue_bits_lo__T_47_mask = 1'h0;
  assign queue_bits_lo__T_47_en = 1'h0;
  assign queue_bits_lo__T_48_data = 32'h0;
  assign queue_bits_lo__T_48_addr = 6'h2b;
  assign queue_bits_lo__T_48_mask = 1'h0;
  assign queue_bits_lo__T_48_en = 1'h0;
  assign queue_bits_lo__T_49_data = 32'h0;
  assign queue_bits_lo__T_49_addr = 6'h2c;
  assign queue_bits_lo__T_49_mask = 1'h0;
  assign queue_bits_lo__T_49_en = 1'h0;
  assign queue_bits_lo__T_50_data = 32'h0;
  assign queue_bits_lo__T_50_addr = 6'h2d;
  assign queue_bits_lo__T_50_mask = 1'h0;
  assign queue_bits_lo__T_50_en = 1'h0;
  assign queue_bits_lo__T_51_data = 32'h0;
  assign queue_bits_lo__T_51_addr = 6'h2e;
  assign queue_bits_lo__T_51_mask = 1'h0;
  assign queue_bits_lo__T_51_en = 1'h0;
  assign queue_bits_lo__T_52_data = 32'h0;
  assign queue_bits_lo__T_52_addr = 6'h2f;
  assign queue_bits_lo__T_52_mask = 1'h0;
  assign queue_bits_lo__T_52_en = 1'h0;
  assign queue_bits_lo__T_53_data = 32'h0;
  assign queue_bits_lo__T_53_addr = 6'h30;
  assign queue_bits_lo__T_53_mask = 1'h0;
  assign queue_bits_lo__T_53_en = 1'h0;
  assign queue_bits_lo__T_54_data = 32'h0;
  assign queue_bits_lo__T_54_addr = 6'h31;
  assign queue_bits_lo__T_54_mask = 1'h0;
  assign queue_bits_lo__T_54_en = 1'h0;
  assign queue_bits_lo__T_55_data = 32'h0;
  assign queue_bits_lo__T_55_addr = 6'h32;
  assign queue_bits_lo__T_55_mask = 1'h0;
  assign queue_bits_lo__T_55_en = 1'h0;
  assign queue_bits_lo__T_56_data = 32'h0;
  assign queue_bits_lo__T_56_addr = 6'h33;
  assign queue_bits_lo__T_56_mask = 1'h0;
  assign queue_bits_lo__T_56_en = 1'h0;
  assign queue_bits_lo__T_57_data = 32'h0;
  assign queue_bits_lo__T_57_addr = 6'h34;
  assign queue_bits_lo__T_57_mask = 1'h0;
  assign queue_bits_lo__T_57_en = 1'h0;
  assign queue_bits_lo__T_58_data = 32'h0;
  assign queue_bits_lo__T_58_addr = 6'h35;
  assign queue_bits_lo__T_58_mask = 1'h0;
  assign queue_bits_lo__T_58_en = 1'h0;
  assign queue_bits_lo__T_59_data = 32'h0;
  assign queue_bits_lo__T_59_addr = 6'h36;
  assign queue_bits_lo__T_59_mask = 1'h0;
  assign queue_bits_lo__T_59_en = 1'h0;
  assign queue_bits_lo__T_60_data = 32'h0;
  assign queue_bits_lo__T_60_addr = 6'h37;
  assign queue_bits_lo__T_60_mask = 1'h0;
  assign queue_bits_lo__T_60_en = 1'h0;
  assign queue_bits_lo__T_61_data = 32'h0;
  assign queue_bits_lo__T_61_addr = 6'h38;
  assign queue_bits_lo__T_61_mask = 1'h0;
  assign queue_bits_lo__T_61_en = 1'h0;
  assign queue_bits_lo__T_62_data = 32'h0;
  assign queue_bits_lo__T_62_addr = 6'h39;
  assign queue_bits_lo__T_62_mask = 1'h0;
  assign queue_bits_lo__T_62_en = 1'h0;
  assign queue_bits_lo__T_63_data = 32'h0;
  assign queue_bits_lo__T_63_addr = 6'h3a;
  assign queue_bits_lo__T_63_mask = 1'h0;
  assign queue_bits_lo__T_63_en = 1'h0;
  assign queue_bits_lo__T_64_data = 32'h0;
  assign queue_bits_lo__T_64_addr = 6'h3b;
  assign queue_bits_lo__T_64_mask = 1'h0;
  assign queue_bits_lo__T_64_en = 1'h0;
  assign queue_bits_lo__T_65_data = 32'h0;
  assign queue_bits_lo__T_65_addr = 6'h3c;
  assign queue_bits_lo__T_65_mask = 1'h0;
  assign queue_bits_lo__T_65_en = 1'h0;
  assign queue_bits_lo__T_66_data = 32'h0;
  assign queue_bits_lo__T_66_addr = 6'h3d;
  assign queue_bits_lo__T_66_mask = 1'h0;
  assign queue_bits_lo__T_66_en = 1'h0;
  assign queue_bits_lo__T_67_data = 32'h0;
  assign queue_bits_lo__T_67_addr = 6'h3e;
  assign queue_bits_lo__T_67_mask = 1'h0;
  assign queue_bits_lo__T_67_en = 1'h0;
  assign queue_bits_lo__T_68_data = 32'h0;
  assign queue_bits_lo__T_68_addr = 6'h3f;
  assign queue_bits_lo__T_68_mask = 1'h0;
  assign queue_bits_lo__T_68_en = 1'h0;
  assign queue_bits_lo__T_70_data = 32'h0;
  assign queue_bits_lo__T_70_addr = 6'h0;
  assign queue_bits_lo__T_70_mask = 1'h0;
  assign queue_bits_lo__T_70_en = reset;
  assign queue_bits_lo__T_71_data = 32'h0;
  assign queue_bits_lo__T_71_addr = 6'h1;
  assign queue_bits_lo__T_71_mask = 1'h0;
  assign queue_bits_lo__T_71_en = reset;
  assign queue_bits_lo__T_72_data = 32'h0;
  assign queue_bits_lo__T_72_addr = 6'h2;
  assign queue_bits_lo__T_72_mask = 1'h0;
  assign queue_bits_lo__T_72_en = reset;
  assign queue_bits_lo__T_73_data = 32'h0;
  assign queue_bits_lo__T_73_addr = 6'h3;
  assign queue_bits_lo__T_73_mask = 1'h0;
  assign queue_bits_lo__T_73_en = reset;
  assign queue_bits_lo__T_74_data = 32'h0;
  assign queue_bits_lo__T_74_addr = 6'h4;
  assign queue_bits_lo__T_74_mask = 1'h0;
  assign queue_bits_lo__T_74_en = reset;
  assign queue_bits_lo__T_75_data = 32'h0;
  assign queue_bits_lo__T_75_addr = 6'h5;
  assign queue_bits_lo__T_75_mask = 1'h0;
  assign queue_bits_lo__T_75_en = reset;
  assign queue_bits_lo__T_76_data = 32'h0;
  assign queue_bits_lo__T_76_addr = 6'h6;
  assign queue_bits_lo__T_76_mask = 1'h0;
  assign queue_bits_lo__T_76_en = reset;
  assign queue_bits_lo__T_77_data = 32'h0;
  assign queue_bits_lo__T_77_addr = 6'h7;
  assign queue_bits_lo__T_77_mask = 1'h0;
  assign queue_bits_lo__T_77_en = reset;
  assign queue_bits_lo__T_78_data = 32'h0;
  assign queue_bits_lo__T_78_addr = 6'h8;
  assign queue_bits_lo__T_78_mask = 1'h0;
  assign queue_bits_lo__T_78_en = reset;
  assign queue_bits_lo__T_79_data = 32'h0;
  assign queue_bits_lo__T_79_addr = 6'h9;
  assign queue_bits_lo__T_79_mask = 1'h0;
  assign queue_bits_lo__T_79_en = reset;
  assign queue_bits_lo__T_80_data = 32'h0;
  assign queue_bits_lo__T_80_addr = 6'ha;
  assign queue_bits_lo__T_80_mask = 1'h0;
  assign queue_bits_lo__T_80_en = reset;
  assign queue_bits_lo__T_81_data = 32'h0;
  assign queue_bits_lo__T_81_addr = 6'hb;
  assign queue_bits_lo__T_81_mask = 1'h0;
  assign queue_bits_lo__T_81_en = reset;
  assign queue_bits_lo__T_82_data = 32'h0;
  assign queue_bits_lo__T_82_addr = 6'hc;
  assign queue_bits_lo__T_82_mask = 1'h0;
  assign queue_bits_lo__T_82_en = reset;
  assign queue_bits_lo__T_83_data = 32'h0;
  assign queue_bits_lo__T_83_addr = 6'hd;
  assign queue_bits_lo__T_83_mask = 1'h0;
  assign queue_bits_lo__T_83_en = reset;
  assign queue_bits_lo__T_84_data = 32'h0;
  assign queue_bits_lo__T_84_addr = 6'he;
  assign queue_bits_lo__T_84_mask = 1'h0;
  assign queue_bits_lo__T_84_en = reset;
  assign queue_bits_lo__T_85_data = 32'h0;
  assign queue_bits_lo__T_85_addr = 6'hf;
  assign queue_bits_lo__T_85_mask = 1'h0;
  assign queue_bits_lo__T_85_en = reset;
  assign queue_bits_lo__T_86_data = 32'h0;
  assign queue_bits_lo__T_86_addr = 6'h10;
  assign queue_bits_lo__T_86_mask = 1'h0;
  assign queue_bits_lo__T_86_en = reset;
  assign queue_bits_lo__T_87_data = 32'h0;
  assign queue_bits_lo__T_87_addr = 6'h11;
  assign queue_bits_lo__T_87_mask = 1'h0;
  assign queue_bits_lo__T_87_en = reset;
  assign queue_bits_lo__T_88_data = 32'h0;
  assign queue_bits_lo__T_88_addr = 6'h12;
  assign queue_bits_lo__T_88_mask = 1'h0;
  assign queue_bits_lo__T_88_en = reset;
  assign queue_bits_lo__T_89_data = 32'h0;
  assign queue_bits_lo__T_89_addr = 6'h13;
  assign queue_bits_lo__T_89_mask = 1'h0;
  assign queue_bits_lo__T_89_en = reset;
  assign queue_bits_lo__T_90_data = 32'h0;
  assign queue_bits_lo__T_90_addr = 6'h14;
  assign queue_bits_lo__T_90_mask = 1'h0;
  assign queue_bits_lo__T_90_en = reset;
  assign queue_bits_lo__T_91_data = 32'h0;
  assign queue_bits_lo__T_91_addr = 6'h15;
  assign queue_bits_lo__T_91_mask = 1'h0;
  assign queue_bits_lo__T_91_en = reset;
  assign queue_bits_lo__T_92_data = 32'h0;
  assign queue_bits_lo__T_92_addr = 6'h16;
  assign queue_bits_lo__T_92_mask = 1'h0;
  assign queue_bits_lo__T_92_en = reset;
  assign queue_bits_lo__T_93_data = 32'h0;
  assign queue_bits_lo__T_93_addr = 6'h17;
  assign queue_bits_lo__T_93_mask = 1'h0;
  assign queue_bits_lo__T_93_en = reset;
  assign queue_bits_lo__T_94_data = 32'h0;
  assign queue_bits_lo__T_94_addr = 6'h18;
  assign queue_bits_lo__T_94_mask = 1'h0;
  assign queue_bits_lo__T_94_en = reset;
  assign queue_bits_lo__T_95_data = 32'h0;
  assign queue_bits_lo__T_95_addr = 6'h19;
  assign queue_bits_lo__T_95_mask = 1'h0;
  assign queue_bits_lo__T_95_en = reset;
  assign queue_bits_lo__T_96_data = 32'h0;
  assign queue_bits_lo__T_96_addr = 6'h1a;
  assign queue_bits_lo__T_96_mask = 1'h0;
  assign queue_bits_lo__T_96_en = reset;
  assign queue_bits_lo__T_97_data = 32'h0;
  assign queue_bits_lo__T_97_addr = 6'h1b;
  assign queue_bits_lo__T_97_mask = 1'h0;
  assign queue_bits_lo__T_97_en = reset;
  assign queue_bits_lo__T_98_data = 32'h0;
  assign queue_bits_lo__T_98_addr = 6'h1c;
  assign queue_bits_lo__T_98_mask = 1'h0;
  assign queue_bits_lo__T_98_en = reset;
  assign queue_bits_lo__T_99_data = 32'h0;
  assign queue_bits_lo__T_99_addr = 6'h1d;
  assign queue_bits_lo__T_99_mask = 1'h0;
  assign queue_bits_lo__T_99_en = reset;
  assign queue_bits_lo__T_100_data = 32'h0;
  assign queue_bits_lo__T_100_addr = 6'h1e;
  assign queue_bits_lo__T_100_mask = 1'h0;
  assign queue_bits_lo__T_100_en = reset;
  assign queue_bits_lo__T_101_data = 32'h0;
  assign queue_bits_lo__T_101_addr = 6'h1f;
  assign queue_bits_lo__T_101_mask = 1'h0;
  assign queue_bits_lo__T_101_en = reset;
  assign queue_bits_lo__T_102_data = 32'h0;
  assign queue_bits_lo__T_102_addr = 6'h20;
  assign queue_bits_lo__T_102_mask = 1'h0;
  assign queue_bits_lo__T_102_en = reset;
  assign queue_bits_lo__T_103_data = 32'h0;
  assign queue_bits_lo__T_103_addr = 6'h21;
  assign queue_bits_lo__T_103_mask = 1'h0;
  assign queue_bits_lo__T_103_en = reset;
  assign queue_bits_lo__T_104_data = 32'h0;
  assign queue_bits_lo__T_104_addr = 6'h22;
  assign queue_bits_lo__T_104_mask = 1'h0;
  assign queue_bits_lo__T_104_en = reset;
  assign queue_bits_lo__T_105_data = 32'h0;
  assign queue_bits_lo__T_105_addr = 6'h23;
  assign queue_bits_lo__T_105_mask = 1'h0;
  assign queue_bits_lo__T_105_en = reset;
  assign queue_bits_lo__T_106_data = 32'h0;
  assign queue_bits_lo__T_106_addr = 6'h24;
  assign queue_bits_lo__T_106_mask = 1'h0;
  assign queue_bits_lo__T_106_en = reset;
  assign queue_bits_lo__T_107_data = 32'h0;
  assign queue_bits_lo__T_107_addr = 6'h25;
  assign queue_bits_lo__T_107_mask = 1'h0;
  assign queue_bits_lo__T_107_en = reset;
  assign queue_bits_lo__T_108_data = 32'h0;
  assign queue_bits_lo__T_108_addr = 6'h26;
  assign queue_bits_lo__T_108_mask = 1'h0;
  assign queue_bits_lo__T_108_en = reset;
  assign queue_bits_lo__T_109_data = 32'h0;
  assign queue_bits_lo__T_109_addr = 6'h27;
  assign queue_bits_lo__T_109_mask = 1'h0;
  assign queue_bits_lo__T_109_en = reset;
  assign queue_bits_lo__T_110_data = 32'h0;
  assign queue_bits_lo__T_110_addr = 6'h28;
  assign queue_bits_lo__T_110_mask = 1'h0;
  assign queue_bits_lo__T_110_en = reset;
  assign queue_bits_lo__T_111_data = 32'h0;
  assign queue_bits_lo__T_111_addr = 6'h29;
  assign queue_bits_lo__T_111_mask = 1'h0;
  assign queue_bits_lo__T_111_en = reset;
  assign queue_bits_lo__T_112_data = 32'h0;
  assign queue_bits_lo__T_112_addr = 6'h2a;
  assign queue_bits_lo__T_112_mask = 1'h0;
  assign queue_bits_lo__T_112_en = reset;
  assign queue_bits_lo__T_113_data = 32'h0;
  assign queue_bits_lo__T_113_addr = 6'h2b;
  assign queue_bits_lo__T_113_mask = 1'h0;
  assign queue_bits_lo__T_113_en = reset;
  assign queue_bits_lo__T_114_data = 32'h0;
  assign queue_bits_lo__T_114_addr = 6'h2c;
  assign queue_bits_lo__T_114_mask = 1'h0;
  assign queue_bits_lo__T_114_en = reset;
  assign queue_bits_lo__T_115_data = 32'h0;
  assign queue_bits_lo__T_115_addr = 6'h2d;
  assign queue_bits_lo__T_115_mask = 1'h0;
  assign queue_bits_lo__T_115_en = reset;
  assign queue_bits_lo__T_116_data = 32'h0;
  assign queue_bits_lo__T_116_addr = 6'h2e;
  assign queue_bits_lo__T_116_mask = 1'h0;
  assign queue_bits_lo__T_116_en = reset;
  assign queue_bits_lo__T_117_data = 32'h0;
  assign queue_bits_lo__T_117_addr = 6'h2f;
  assign queue_bits_lo__T_117_mask = 1'h0;
  assign queue_bits_lo__T_117_en = reset;
  assign queue_bits_lo__T_118_data = 32'h0;
  assign queue_bits_lo__T_118_addr = 6'h30;
  assign queue_bits_lo__T_118_mask = 1'h0;
  assign queue_bits_lo__T_118_en = reset;
  assign queue_bits_lo__T_119_data = 32'h0;
  assign queue_bits_lo__T_119_addr = 6'h31;
  assign queue_bits_lo__T_119_mask = 1'h0;
  assign queue_bits_lo__T_119_en = reset;
  assign queue_bits_lo__T_120_data = 32'h0;
  assign queue_bits_lo__T_120_addr = 6'h32;
  assign queue_bits_lo__T_120_mask = 1'h0;
  assign queue_bits_lo__T_120_en = reset;
  assign queue_bits_lo__T_121_data = 32'h0;
  assign queue_bits_lo__T_121_addr = 6'h33;
  assign queue_bits_lo__T_121_mask = 1'h0;
  assign queue_bits_lo__T_121_en = reset;
  assign queue_bits_lo__T_122_data = 32'h0;
  assign queue_bits_lo__T_122_addr = 6'h34;
  assign queue_bits_lo__T_122_mask = 1'h0;
  assign queue_bits_lo__T_122_en = reset;
  assign queue_bits_lo__T_123_data = 32'h0;
  assign queue_bits_lo__T_123_addr = 6'h35;
  assign queue_bits_lo__T_123_mask = 1'h0;
  assign queue_bits_lo__T_123_en = reset;
  assign queue_bits_lo__T_124_data = 32'h0;
  assign queue_bits_lo__T_124_addr = 6'h36;
  assign queue_bits_lo__T_124_mask = 1'h0;
  assign queue_bits_lo__T_124_en = reset;
  assign queue_bits_lo__T_125_data = 32'h0;
  assign queue_bits_lo__T_125_addr = 6'h37;
  assign queue_bits_lo__T_125_mask = 1'h0;
  assign queue_bits_lo__T_125_en = reset;
  assign queue_bits_lo__T_126_data = 32'h0;
  assign queue_bits_lo__T_126_addr = 6'h38;
  assign queue_bits_lo__T_126_mask = 1'h0;
  assign queue_bits_lo__T_126_en = reset;
  assign queue_bits_lo__T_127_data = 32'h0;
  assign queue_bits_lo__T_127_addr = 6'h39;
  assign queue_bits_lo__T_127_mask = 1'h0;
  assign queue_bits_lo__T_127_en = reset;
  assign queue_bits_lo__T_128_data = 32'h0;
  assign queue_bits_lo__T_128_addr = 6'h3a;
  assign queue_bits_lo__T_128_mask = 1'h0;
  assign queue_bits_lo__T_128_en = reset;
  assign queue_bits_lo__T_129_data = 32'h0;
  assign queue_bits_lo__T_129_addr = 6'h3b;
  assign queue_bits_lo__T_129_mask = 1'h0;
  assign queue_bits_lo__T_129_en = reset;
  assign queue_bits_lo__T_130_data = 32'h0;
  assign queue_bits_lo__T_130_addr = 6'h3c;
  assign queue_bits_lo__T_130_mask = 1'h0;
  assign queue_bits_lo__T_130_en = reset;
  assign queue_bits_lo__T_131_data = 32'h0;
  assign queue_bits_lo__T_131_addr = 6'h3d;
  assign queue_bits_lo__T_131_mask = 1'h0;
  assign queue_bits_lo__T_131_en = reset;
  assign queue_bits_lo__T_132_data = 32'h0;
  assign queue_bits_lo__T_132_addr = 6'h3e;
  assign queue_bits_lo__T_132_mask = 1'h0;
  assign queue_bits_lo__T_132_en = reset;
  assign queue_bits_lo__T_133_data = 32'h0;
  assign queue_bits_lo__T_133_addr = 6'h3f;
  assign queue_bits_lo__T_133_mask = 1'h0;
  assign queue_bits_lo__T_133_en = reset;
  assign queue_bits_lo_q_head_w_data = 32'h0;
  assign queue_bits_lo_q_head_w_addr = head;
  assign queue_bits_lo_q_head_w_mask = 1'h0;
  assign queue_bits_lo_q_head_w_en = io_deq_valid;
  assign queue_bits_op1_q_head_r_addr = head;
  assign queue_bits_op1_q_head_r_data = queue_bits_op1[queue_bits_op1_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_op1__T_3_data = io_enq_0_bits_data_op1;
  assign queue_bits_op1__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_op1__T_3_mask = 1'h1;
  assign queue_bits_op1__T_3_en = io_enq_0_valid;
  assign queue_bits_op1__T_4_data = io_enq_1_bits_data_op1;
  assign queue_bits_op1__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_op1__T_4_mask = 1'h1;
  assign queue_bits_op1__T_4_en = io_enq_1_valid;
  assign queue_bits_op1__T_5_data = 32'h0;
  assign queue_bits_op1__T_5_addr = 6'h0;
  assign queue_bits_op1__T_5_mask = 1'h0;
  assign queue_bits_op1__T_5_en = 1'h0;
  assign queue_bits_op1__T_6_data = 32'h0;
  assign queue_bits_op1__T_6_addr = 6'h1;
  assign queue_bits_op1__T_6_mask = 1'h0;
  assign queue_bits_op1__T_6_en = 1'h0;
  assign queue_bits_op1__T_7_data = 32'h0;
  assign queue_bits_op1__T_7_addr = 6'h2;
  assign queue_bits_op1__T_7_mask = 1'h0;
  assign queue_bits_op1__T_7_en = 1'h0;
  assign queue_bits_op1__T_8_data = 32'h0;
  assign queue_bits_op1__T_8_addr = 6'h3;
  assign queue_bits_op1__T_8_mask = 1'h0;
  assign queue_bits_op1__T_8_en = 1'h0;
  assign queue_bits_op1__T_9_data = 32'h0;
  assign queue_bits_op1__T_9_addr = 6'h4;
  assign queue_bits_op1__T_9_mask = 1'h0;
  assign queue_bits_op1__T_9_en = 1'h0;
  assign queue_bits_op1__T_10_data = 32'h0;
  assign queue_bits_op1__T_10_addr = 6'h5;
  assign queue_bits_op1__T_10_mask = 1'h0;
  assign queue_bits_op1__T_10_en = 1'h0;
  assign queue_bits_op1__T_11_data = 32'h0;
  assign queue_bits_op1__T_11_addr = 6'h6;
  assign queue_bits_op1__T_11_mask = 1'h0;
  assign queue_bits_op1__T_11_en = 1'h0;
  assign queue_bits_op1__T_12_data = 32'h0;
  assign queue_bits_op1__T_12_addr = 6'h7;
  assign queue_bits_op1__T_12_mask = 1'h0;
  assign queue_bits_op1__T_12_en = 1'h0;
  assign queue_bits_op1__T_13_data = 32'h0;
  assign queue_bits_op1__T_13_addr = 6'h8;
  assign queue_bits_op1__T_13_mask = 1'h0;
  assign queue_bits_op1__T_13_en = 1'h0;
  assign queue_bits_op1__T_14_data = 32'h0;
  assign queue_bits_op1__T_14_addr = 6'h9;
  assign queue_bits_op1__T_14_mask = 1'h0;
  assign queue_bits_op1__T_14_en = 1'h0;
  assign queue_bits_op1__T_15_data = 32'h0;
  assign queue_bits_op1__T_15_addr = 6'ha;
  assign queue_bits_op1__T_15_mask = 1'h0;
  assign queue_bits_op1__T_15_en = 1'h0;
  assign queue_bits_op1__T_16_data = 32'h0;
  assign queue_bits_op1__T_16_addr = 6'hb;
  assign queue_bits_op1__T_16_mask = 1'h0;
  assign queue_bits_op1__T_16_en = 1'h0;
  assign queue_bits_op1__T_17_data = 32'h0;
  assign queue_bits_op1__T_17_addr = 6'hc;
  assign queue_bits_op1__T_17_mask = 1'h0;
  assign queue_bits_op1__T_17_en = 1'h0;
  assign queue_bits_op1__T_18_data = 32'h0;
  assign queue_bits_op1__T_18_addr = 6'hd;
  assign queue_bits_op1__T_18_mask = 1'h0;
  assign queue_bits_op1__T_18_en = 1'h0;
  assign queue_bits_op1__T_19_data = 32'h0;
  assign queue_bits_op1__T_19_addr = 6'he;
  assign queue_bits_op1__T_19_mask = 1'h0;
  assign queue_bits_op1__T_19_en = 1'h0;
  assign queue_bits_op1__T_20_data = 32'h0;
  assign queue_bits_op1__T_20_addr = 6'hf;
  assign queue_bits_op1__T_20_mask = 1'h0;
  assign queue_bits_op1__T_20_en = 1'h0;
  assign queue_bits_op1__T_21_data = 32'h0;
  assign queue_bits_op1__T_21_addr = 6'h10;
  assign queue_bits_op1__T_21_mask = 1'h0;
  assign queue_bits_op1__T_21_en = 1'h0;
  assign queue_bits_op1__T_22_data = 32'h0;
  assign queue_bits_op1__T_22_addr = 6'h11;
  assign queue_bits_op1__T_22_mask = 1'h0;
  assign queue_bits_op1__T_22_en = 1'h0;
  assign queue_bits_op1__T_23_data = 32'h0;
  assign queue_bits_op1__T_23_addr = 6'h12;
  assign queue_bits_op1__T_23_mask = 1'h0;
  assign queue_bits_op1__T_23_en = 1'h0;
  assign queue_bits_op1__T_24_data = 32'h0;
  assign queue_bits_op1__T_24_addr = 6'h13;
  assign queue_bits_op1__T_24_mask = 1'h0;
  assign queue_bits_op1__T_24_en = 1'h0;
  assign queue_bits_op1__T_25_data = 32'h0;
  assign queue_bits_op1__T_25_addr = 6'h14;
  assign queue_bits_op1__T_25_mask = 1'h0;
  assign queue_bits_op1__T_25_en = 1'h0;
  assign queue_bits_op1__T_26_data = 32'h0;
  assign queue_bits_op1__T_26_addr = 6'h15;
  assign queue_bits_op1__T_26_mask = 1'h0;
  assign queue_bits_op1__T_26_en = 1'h0;
  assign queue_bits_op1__T_27_data = 32'h0;
  assign queue_bits_op1__T_27_addr = 6'h16;
  assign queue_bits_op1__T_27_mask = 1'h0;
  assign queue_bits_op1__T_27_en = 1'h0;
  assign queue_bits_op1__T_28_data = 32'h0;
  assign queue_bits_op1__T_28_addr = 6'h17;
  assign queue_bits_op1__T_28_mask = 1'h0;
  assign queue_bits_op1__T_28_en = 1'h0;
  assign queue_bits_op1__T_29_data = 32'h0;
  assign queue_bits_op1__T_29_addr = 6'h18;
  assign queue_bits_op1__T_29_mask = 1'h0;
  assign queue_bits_op1__T_29_en = 1'h0;
  assign queue_bits_op1__T_30_data = 32'h0;
  assign queue_bits_op1__T_30_addr = 6'h19;
  assign queue_bits_op1__T_30_mask = 1'h0;
  assign queue_bits_op1__T_30_en = 1'h0;
  assign queue_bits_op1__T_31_data = 32'h0;
  assign queue_bits_op1__T_31_addr = 6'h1a;
  assign queue_bits_op1__T_31_mask = 1'h0;
  assign queue_bits_op1__T_31_en = 1'h0;
  assign queue_bits_op1__T_32_data = 32'h0;
  assign queue_bits_op1__T_32_addr = 6'h1b;
  assign queue_bits_op1__T_32_mask = 1'h0;
  assign queue_bits_op1__T_32_en = 1'h0;
  assign queue_bits_op1__T_33_data = 32'h0;
  assign queue_bits_op1__T_33_addr = 6'h1c;
  assign queue_bits_op1__T_33_mask = 1'h0;
  assign queue_bits_op1__T_33_en = 1'h0;
  assign queue_bits_op1__T_34_data = 32'h0;
  assign queue_bits_op1__T_34_addr = 6'h1d;
  assign queue_bits_op1__T_34_mask = 1'h0;
  assign queue_bits_op1__T_34_en = 1'h0;
  assign queue_bits_op1__T_35_data = 32'h0;
  assign queue_bits_op1__T_35_addr = 6'h1e;
  assign queue_bits_op1__T_35_mask = 1'h0;
  assign queue_bits_op1__T_35_en = 1'h0;
  assign queue_bits_op1__T_36_data = 32'h0;
  assign queue_bits_op1__T_36_addr = 6'h1f;
  assign queue_bits_op1__T_36_mask = 1'h0;
  assign queue_bits_op1__T_36_en = 1'h0;
  assign queue_bits_op1__T_37_data = 32'h0;
  assign queue_bits_op1__T_37_addr = 6'h20;
  assign queue_bits_op1__T_37_mask = 1'h0;
  assign queue_bits_op1__T_37_en = 1'h0;
  assign queue_bits_op1__T_38_data = 32'h0;
  assign queue_bits_op1__T_38_addr = 6'h21;
  assign queue_bits_op1__T_38_mask = 1'h0;
  assign queue_bits_op1__T_38_en = 1'h0;
  assign queue_bits_op1__T_39_data = 32'h0;
  assign queue_bits_op1__T_39_addr = 6'h22;
  assign queue_bits_op1__T_39_mask = 1'h0;
  assign queue_bits_op1__T_39_en = 1'h0;
  assign queue_bits_op1__T_40_data = 32'h0;
  assign queue_bits_op1__T_40_addr = 6'h23;
  assign queue_bits_op1__T_40_mask = 1'h0;
  assign queue_bits_op1__T_40_en = 1'h0;
  assign queue_bits_op1__T_41_data = 32'h0;
  assign queue_bits_op1__T_41_addr = 6'h24;
  assign queue_bits_op1__T_41_mask = 1'h0;
  assign queue_bits_op1__T_41_en = 1'h0;
  assign queue_bits_op1__T_42_data = 32'h0;
  assign queue_bits_op1__T_42_addr = 6'h25;
  assign queue_bits_op1__T_42_mask = 1'h0;
  assign queue_bits_op1__T_42_en = 1'h0;
  assign queue_bits_op1__T_43_data = 32'h0;
  assign queue_bits_op1__T_43_addr = 6'h26;
  assign queue_bits_op1__T_43_mask = 1'h0;
  assign queue_bits_op1__T_43_en = 1'h0;
  assign queue_bits_op1__T_44_data = 32'h0;
  assign queue_bits_op1__T_44_addr = 6'h27;
  assign queue_bits_op1__T_44_mask = 1'h0;
  assign queue_bits_op1__T_44_en = 1'h0;
  assign queue_bits_op1__T_45_data = 32'h0;
  assign queue_bits_op1__T_45_addr = 6'h28;
  assign queue_bits_op1__T_45_mask = 1'h0;
  assign queue_bits_op1__T_45_en = 1'h0;
  assign queue_bits_op1__T_46_data = 32'h0;
  assign queue_bits_op1__T_46_addr = 6'h29;
  assign queue_bits_op1__T_46_mask = 1'h0;
  assign queue_bits_op1__T_46_en = 1'h0;
  assign queue_bits_op1__T_47_data = 32'h0;
  assign queue_bits_op1__T_47_addr = 6'h2a;
  assign queue_bits_op1__T_47_mask = 1'h0;
  assign queue_bits_op1__T_47_en = 1'h0;
  assign queue_bits_op1__T_48_data = 32'h0;
  assign queue_bits_op1__T_48_addr = 6'h2b;
  assign queue_bits_op1__T_48_mask = 1'h0;
  assign queue_bits_op1__T_48_en = 1'h0;
  assign queue_bits_op1__T_49_data = 32'h0;
  assign queue_bits_op1__T_49_addr = 6'h2c;
  assign queue_bits_op1__T_49_mask = 1'h0;
  assign queue_bits_op1__T_49_en = 1'h0;
  assign queue_bits_op1__T_50_data = 32'h0;
  assign queue_bits_op1__T_50_addr = 6'h2d;
  assign queue_bits_op1__T_50_mask = 1'h0;
  assign queue_bits_op1__T_50_en = 1'h0;
  assign queue_bits_op1__T_51_data = 32'h0;
  assign queue_bits_op1__T_51_addr = 6'h2e;
  assign queue_bits_op1__T_51_mask = 1'h0;
  assign queue_bits_op1__T_51_en = 1'h0;
  assign queue_bits_op1__T_52_data = 32'h0;
  assign queue_bits_op1__T_52_addr = 6'h2f;
  assign queue_bits_op1__T_52_mask = 1'h0;
  assign queue_bits_op1__T_52_en = 1'h0;
  assign queue_bits_op1__T_53_data = 32'h0;
  assign queue_bits_op1__T_53_addr = 6'h30;
  assign queue_bits_op1__T_53_mask = 1'h0;
  assign queue_bits_op1__T_53_en = 1'h0;
  assign queue_bits_op1__T_54_data = 32'h0;
  assign queue_bits_op1__T_54_addr = 6'h31;
  assign queue_bits_op1__T_54_mask = 1'h0;
  assign queue_bits_op1__T_54_en = 1'h0;
  assign queue_bits_op1__T_55_data = 32'h0;
  assign queue_bits_op1__T_55_addr = 6'h32;
  assign queue_bits_op1__T_55_mask = 1'h0;
  assign queue_bits_op1__T_55_en = 1'h0;
  assign queue_bits_op1__T_56_data = 32'h0;
  assign queue_bits_op1__T_56_addr = 6'h33;
  assign queue_bits_op1__T_56_mask = 1'h0;
  assign queue_bits_op1__T_56_en = 1'h0;
  assign queue_bits_op1__T_57_data = 32'h0;
  assign queue_bits_op1__T_57_addr = 6'h34;
  assign queue_bits_op1__T_57_mask = 1'h0;
  assign queue_bits_op1__T_57_en = 1'h0;
  assign queue_bits_op1__T_58_data = 32'h0;
  assign queue_bits_op1__T_58_addr = 6'h35;
  assign queue_bits_op1__T_58_mask = 1'h0;
  assign queue_bits_op1__T_58_en = 1'h0;
  assign queue_bits_op1__T_59_data = 32'h0;
  assign queue_bits_op1__T_59_addr = 6'h36;
  assign queue_bits_op1__T_59_mask = 1'h0;
  assign queue_bits_op1__T_59_en = 1'h0;
  assign queue_bits_op1__T_60_data = 32'h0;
  assign queue_bits_op1__T_60_addr = 6'h37;
  assign queue_bits_op1__T_60_mask = 1'h0;
  assign queue_bits_op1__T_60_en = 1'h0;
  assign queue_bits_op1__T_61_data = 32'h0;
  assign queue_bits_op1__T_61_addr = 6'h38;
  assign queue_bits_op1__T_61_mask = 1'h0;
  assign queue_bits_op1__T_61_en = 1'h0;
  assign queue_bits_op1__T_62_data = 32'h0;
  assign queue_bits_op1__T_62_addr = 6'h39;
  assign queue_bits_op1__T_62_mask = 1'h0;
  assign queue_bits_op1__T_62_en = 1'h0;
  assign queue_bits_op1__T_63_data = 32'h0;
  assign queue_bits_op1__T_63_addr = 6'h3a;
  assign queue_bits_op1__T_63_mask = 1'h0;
  assign queue_bits_op1__T_63_en = 1'h0;
  assign queue_bits_op1__T_64_data = 32'h0;
  assign queue_bits_op1__T_64_addr = 6'h3b;
  assign queue_bits_op1__T_64_mask = 1'h0;
  assign queue_bits_op1__T_64_en = 1'h0;
  assign queue_bits_op1__T_65_data = 32'h0;
  assign queue_bits_op1__T_65_addr = 6'h3c;
  assign queue_bits_op1__T_65_mask = 1'h0;
  assign queue_bits_op1__T_65_en = 1'h0;
  assign queue_bits_op1__T_66_data = 32'h0;
  assign queue_bits_op1__T_66_addr = 6'h3d;
  assign queue_bits_op1__T_66_mask = 1'h0;
  assign queue_bits_op1__T_66_en = 1'h0;
  assign queue_bits_op1__T_67_data = 32'h0;
  assign queue_bits_op1__T_67_addr = 6'h3e;
  assign queue_bits_op1__T_67_mask = 1'h0;
  assign queue_bits_op1__T_67_en = 1'h0;
  assign queue_bits_op1__T_68_data = 32'h0;
  assign queue_bits_op1__T_68_addr = 6'h3f;
  assign queue_bits_op1__T_68_mask = 1'h0;
  assign queue_bits_op1__T_68_en = 1'h0;
  assign queue_bits_op1__T_70_data = 32'h0;
  assign queue_bits_op1__T_70_addr = 6'h0;
  assign queue_bits_op1__T_70_mask = 1'h0;
  assign queue_bits_op1__T_70_en = reset;
  assign queue_bits_op1__T_71_data = 32'h0;
  assign queue_bits_op1__T_71_addr = 6'h1;
  assign queue_bits_op1__T_71_mask = 1'h0;
  assign queue_bits_op1__T_71_en = reset;
  assign queue_bits_op1__T_72_data = 32'h0;
  assign queue_bits_op1__T_72_addr = 6'h2;
  assign queue_bits_op1__T_72_mask = 1'h0;
  assign queue_bits_op1__T_72_en = reset;
  assign queue_bits_op1__T_73_data = 32'h0;
  assign queue_bits_op1__T_73_addr = 6'h3;
  assign queue_bits_op1__T_73_mask = 1'h0;
  assign queue_bits_op1__T_73_en = reset;
  assign queue_bits_op1__T_74_data = 32'h0;
  assign queue_bits_op1__T_74_addr = 6'h4;
  assign queue_bits_op1__T_74_mask = 1'h0;
  assign queue_bits_op1__T_74_en = reset;
  assign queue_bits_op1__T_75_data = 32'h0;
  assign queue_bits_op1__T_75_addr = 6'h5;
  assign queue_bits_op1__T_75_mask = 1'h0;
  assign queue_bits_op1__T_75_en = reset;
  assign queue_bits_op1__T_76_data = 32'h0;
  assign queue_bits_op1__T_76_addr = 6'h6;
  assign queue_bits_op1__T_76_mask = 1'h0;
  assign queue_bits_op1__T_76_en = reset;
  assign queue_bits_op1__T_77_data = 32'h0;
  assign queue_bits_op1__T_77_addr = 6'h7;
  assign queue_bits_op1__T_77_mask = 1'h0;
  assign queue_bits_op1__T_77_en = reset;
  assign queue_bits_op1__T_78_data = 32'h0;
  assign queue_bits_op1__T_78_addr = 6'h8;
  assign queue_bits_op1__T_78_mask = 1'h0;
  assign queue_bits_op1__T_78_en = reset;
  assign queue_bits_op1__T_79_data = 32'h0;
  assign queue_bits_op1__T_79_addr = 6'h9;
  assign queue_bits_op1__T_79_mask = 1'h0;
  assign queue_bits_op1__T_79_en = reset;
  assign queue_bits_op1__T_80_data = 32'h0;
  assign queue_bits_op1__T_80_addr = 6'ha;
  assign queue_bits_op1__T_80_mask = 1'h0;
  assign queue_bits_op1__T_80_en = reset;
  assign queue_bits_op1__T_81_data = 32'h0;
  assign queue_bits_op1__T_81_addr = 6'hb;
  assign queue_bits_op1__T_81_mask = 1'h0;
  assign queue_bits_op1__T_81_en = reset;
  assign queue_bits_op1__T_82_data = 32'h0;
  assign queue_bits_op1__T_82_addr = 6'hc;
  assign queue_bits_op1__T_82_mask = 1'h0;
  assign queue_bits_op1__T_82_en = reset;
  assign queue_bits_op1__T_83_data = 32'h0;
  assign queue_bits_op1__T_83_addr = 6'hd;
  assign queue_bits_op1__T_83_mask = 1'h0;
  assign queue_bits_op1__T_83_en = reset;
  assign queue_bits_op1__T_84_data = 32'h0;
  assign queue_bits_op1__T_84_addr = 6'he;
  assign queue_bits_op1__T_84_mask = 1'h0;
  assign queue_bits_op1__T_84_en = reset;
  assign queue_bits_op1__T_85_data = 32'h0;
  assign queue_bits_op1__T_85_addr = 6'hf;
  assign queue_bits_op1__T_85_mask = 1'h0;
  assign queue_bits_op1__T_85_en = reset;
  assign queue_bits_op1__T_86_data = 32'h0;
  assign queue_bits_op1__T_86_addr = 6'h10;
  assign queue_bits_op1__T_86_mask = 1'h0;
  assign queue_bits_op1__T_86_en = reset;
  assign queue_bits_op1__T_87_data = 32'h0;
  assign queue_bits_op1__T_87_addr = 6'h11;
  assign queue_bits_op1__T_87_mask = 1'h0;
  assign queue_bits_op1__T_87_en = reset;
  assign queue_bits_op1__T_88_data = 32'h0;
  assign queue_bits_op1__T_88_addr = 6'h12;
  assign queue_bits_op1__T_88_mask = 1'h0;
  assign queue_bits_op1__T_88_en = reset;
  assign queue_bits_op1__T_89_data = 32'h0;
  assign queue_bits_op1__T_89_addr = 6'h13;
  assign queue_bits_op1__T_89_mask = 1'h0;
  assign queue_bits_op1__T_89_en = reset;
  assign queue_bits_op1__T_90_data = 32'h0;
  assign queue_bits_op1__T_90_addr = 6'h14;
  assign queue_bits_op1__T_90_mask = 1'h0;
  assign queue_bits_op1__T_90_en = reset;
  assign queue_bits_op1__T_91_data = 32'h0;
  assign queue_bits_op1__T_91_addr = 6'h15;
  assign queue_bits_op1__T_91_mask = 1'h0;
  assign queue_bits_op1__T_91_en = reset;
  assign queue_bits_op1__T_92_data = 32'h0;
  assign queue_bits_op1__T_92_addr = 6'h16;
  assign queue_bits_op1__T_92_mask = 1'h0;
  assign queue_bits_op1__T_92_en = reset;
  assign queue_bits_op1__T_93_data = 32'h0;
  assign queue_bits_op1__T_93_addr = 6'h17;
  assign queue_bits_op1__T_93_mask = 1'h0;
  assign queue_bits_op1__T_93_en = reset;
  assign queue_bits_op1__T_94_data = 32'h0;
  assign queue_bits_op1__T_94_addr = 6'h18;
  assign queue_bits_op1__T_94_mask = 1'h0;
  assign queue_bits_op1__T_94_en = reset;
  assign queue_bits_op1__T_95_data = 32'h0;
  assign queue_bits_op1__T_95_addr = 6'h19;
  assign queue_bits_op1__T_95_mask = 1'h0;
  assign queue_bits_op1__T_95_en = reset;
  assign queue_bits_op1__T_96_data = 32'h0;
  assign queue_bits_op1__T_96_addr = 6'h1a;
  assign queue_bits_op1__T_96_mask = 1'h0;
  assign queue_bits_op1__T_96_en = reset;
  assign queue_bits_op1__T_97_data = 32'h0;
  assign queue_bits_op1__T_97_addr = 6'h1b;
  assign queue_bits_op1__T_97_mask = 1'h0;
  assign queue_bits_op1__T_97_en = reset;
  assign queue_bits_op1__T_98_data = 32'h0;
  assign queue_bits_op1__T_98_addr = 6'h1c;
  assign queue_bits_op1__T_98_mask = 1'h0;
  assign queue_bits_op1__T_98_en = reset;
  assign queue_bits_op1__T_99_data = 32'h0;
  assign queue_bits_op1__T_99_addr = 6'h1d;
  assign queue_bits_op1__T_99_mask = 1'h0;
  assign queue_bits_op1__T_99_en = reset;
  assign queue_bits_op1__T_100_data = 32'h0;
  assign queue_bits_op1__T_100_addr = 6'h1e;
  assign queue_bits_op1__T_100_mask = 1'h0;
  assign queue_bits_op1__T_100_en = reset;
  assign queue_bits_op1__T_101_data = 32'h0;
  assign queue_bits_op1__T_101_addr = 6'h1f;
  assign queue_bits_op1__T_101_mask = 1'h0;
  assign queue_bits_op1__T_101_en = reset;
  assign queue_bits_op1__T_102_data = 32'h0;
  assign queue_bits_op1__T_102_addr = 6'h20;
  assign queue_bits_op1__T_102_mask = 1'h0;
  assign queue_bits_op1__T_102_en = reset;
  assign queue_bits_op1__T_103_data = 32'h0;
  assign queue_bits_op1__T_103_addr = 6'h21;
  assign queue_bits_op1__T_103_mask = 1'h0;
  assign queue_bits_op1__T_103_en = reset;
  assign queue_bits_op1__T_104_data = 32'h0;
  assign queue_bits_op1__T_104_addr = 6'h22;
  assign queue_bits_op1__T_104_mask = 1'h0;
  assign queue_bits_op1__T_104_en = reset;
  assign queue_bits_op1__T_105_data = 32'h0;
  assign queue_bits_op1__T_105_addr = 6'h23;
  assign queue_bits_op1__T_105_mask = 1'h0;
  assign queue_bits_op1__T_105_en = reset;
  assign queue_bits_op1__T_106_data = 32'h0;
  assign queue_bits_op1__T_106_addr = 6'h24;
  assign queue_bits_op1__T_106_mask = 1'h0;
  assign queue_bits_op1__T_106_en = reset;
  assign queue_bits_op1__T_107_data = 32'h0;
  assign queue_bits_op1__T_107_addr = 6'h25;
  assign queue_bits_op1__T_107_mask = 1'h0;
  assign queue_bits_op1__T_107_en = reset;
  assign queue_bits_op1__T_108_data = 32'h0;
  assign queue_bits_op1__T_108_addr = 6'h26;
  assign queue_bits_op1__T_108_mask = 1'h0;
  assign queue_bits_op1__T_108_en = reset;
  assign queue_bits_op1__T_109_data = 32'h0;
  assign queue_bits_op1__T_109_addr = 6'h27;
  assign queue_bits_op1__T_109_mask = 1'h0;
  assign queue_bits_op1__T_109_en = reset;
  assign queue_bits_op1__T_110_data = 32'h0;
  assign queue_bits_op1__T_110_addr = 6'h28;
  assign queue_bits_op1__T_110_mask = 1'h0;
  assign queue_bits_op1__T_110_en = reset;
  assign queue_bits_op1__T_111_data = 32'h0;
  assign queue_bits_op1__T_111_addr = 6'h29;
  assign queue_bits_op1__T_111_mask = 1'h0;
  assign queue_bits_op1__T_111_en = reset;
  assign queue_bits_op1__T_112_data = 32'h0;
  assign queue_bits_op1__T_112_addr = 6'h2a;
  assign queue_bits_op1__T_112_mask = 1'h0;
  assign queue_bits_op1__T_112_en = reset;
  assign queue_bits_op1__T_113_data = 32'h0;
  assign queue_bits_op1__T_113_addr = 6'h2b;
  assign queue_bits_op1__T_113_mask = 1'h0;
  assign queue_bits_op1__T_113_en = reset;
  assign queue_bits_op1__T_114_data = 32'h0;
  assign queue_bits_op1__T_114_addr = 6'h2c;
  assign queue_bits_op1__T_114_mask = 1'h0;
  assign queue_bits_op1__T_114_en = reset;
  assign queue_bits_op1__T_115_data = 32'h0;
  assign queue_bits_op1__T_115_addr = 6'h2d;
  assign queue_bits_op1__T_115_mask = 1'h0;
  assign queue_bits_op1__T_115_en = reset;
  assign queue_bits_op1__T_116_data = 32'h0;
  assign queue_bits_op1__T_116_addr = 6'h2e;
  assign queue_bits_op1__T_116_mask = 1'h0;
  assign queue_bits_op1__T_116_en = reset;
  assign queue_bits_op1__T_117_data = 32'h0;
  assign queue_bits_op1__T_117_addr = 6'h2f;
  assign queue_bits_op1__T_117_mask = 1'h0;
  assign queue_bits_op1__T_117_en = reset;
  assign queue_bits_op1__T_118_data = 32'h0;
  assign queue_bits_op1__T_118_addr = 6'h30;
  assign queue_bits_op1__T_118_mask = 1'h0;
  assign queue_bits_op1__T_118_en = reset;
  assign queue_bits_op1__T_119_data = 32'h0;
  assign queue_bits_op1__T_119_addr = 6'h31;
  assign queue_bits_op1__T_119_mask = 1'h0;
  assign queue_bits_op1__T_119_en = reset;
  assign queue_bits_op1__T_120_data = 32'h0;
  assign queue_bits_op1__T_120_addr = 6'h32;
  assign queue_bits_op1__T_120_mask = 1'h0;
  assign queue_bits_op1__T_120_en = reset;
  assign queue_bits_op1__T_121_data = 32'h0;
  assign queue_bits_op1__T_121_addr = 6'h33;
  assign queue_bits_op1__T_121_mask = 1'h0;
  assign queue_bits_op1__T_121_en = reset;
  assign queue_bits_op1__T_122_data = 32'h0;
  assign queue_bits_op1__T_122_addr = 6'h34;
  assign queue_bits_op1__T_122_mask = 1'h0;
  assign queue_bits_op1__T_122_en = reset;
  assign queue_bits_op1__T_123_data = 32'h0;
  assign queue_bits_op1__T_123_addr = 6'h35;
  assign queue_bits_op1__T_123_mask = 1'h0;
  assign queue_bits_op1__T_123_en = reset;
  assign queue_bits_op1__T_124_data = 32'h0;
  assign queue_bits_op1__T_124_addr = 6'h36;
  assign queue_bits_op1__T_124_mask = 1'h0;
  assign queue_bits_op1__T_124_en = reset;
  assign queue_bits_op1__T_125_data = 32'h0;
  assign queue_bits_op1__T_125_addr = 6'h37;
  assign queue_bits_op1__T_125_mask = 1'h0;
  assign queue_bits_op1__T_125_en = reset;
  assign queue_bits_op1__T_126_data = 32'h0;
  assign queue_bits_op1__T_126_addr = 6'h38;
  assign queue_bits_op1__T_126_mask = 1'h0;
  assign queue_bits_op1__T_126_en = reset;
  assign queue_bits_op1__T_127_data = 32'h0;
  assign queue_bits_op1__T_127_addr = 6'h39;
  assign queue_bits_op1__T_127_mask = 1'h0;
  assign queue_bits_op1__T_127_en = reset;
  assign queue_bits_op1__T_128_data = 32'h0;
  assign queue_bits_op1__T_128_addr = 6'h3a;
  assign queue_bits_op1__T_128_mask = 1'h0;
  assign queue_bits_op1__T_128_en = reset;
  assign queue_bits_op1__T_129_data = 32'h0;
  assign queue_bits_op1__T_129_addr = 6'h3b;
  assign queue_bits_op1__T_129_mask = 1'h0;
  assign queue_bits_op1__T_129_en = reset;
  assign queue_bits_op1__T_130_data = 32'h0;
  assign queue_bits_op1__T_130_addr = 6'h3c;
  assign queue_bits_op1__T_130_mask = 1'h0;
  assign queue_bits_op1__T_130_en = reset;
  assign queue_bits_op1__T_131_data = 32'h0;
  assign queue_bits_op1__T_131_addr = 6'h3d;
  assign queue_bits_op1__T_131_mask = 1'h0;
  assign queue_bits_op1__T_131_en = reset;
  assign queue_bits_op1__T_132_data = 32'h0;
  assign queue_bits_op1__T_132_addr = 6'h3e;
  assign queue_bits_op1__T_132_mask = 1'h0;
  assign queue_bits_op1__T_132_en = reset;
  assign queue_bits_op1__T_133_data = 32'h0;
  assign queue_bits_op1__T_133_addr = 6'h3f;
  assign queue_bits_op1__T_133_mask = 1'h0;
  assign queue_bits_op1__T_133_en = reset;
  assign queue_bits_op1_q_head_w_data = 32'h0;
  assign queue_bits_op1_q_head_w_addr = head;
  assign queue_bits_op1_q_head_w_mask = 1'h0;
  assign queue_bits_op1_q_head_w_en = io_deq_valid;
  assign queue_bits_fu_op_q_head_r_addr = head;
  assign queue_bits_fu_op_q_head_r_data = queue_bits_fu_op[queue_bits_fu_op_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_fu_op__T_3_data = io_enq_0_bits_data_fu_op;
  assign queue_bits_fu_op__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_fu_op__T_3_mask = 1'h1;
  assign queue_bits_fu_op__T_3_en = io_enq_0_valid;
  assign queue_bits_fu_op__T_4_data = io_enq_1_bits_data_fu_op;
  assign queue_bits_fu_op__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_fu_op__T_4_mask = 1'h1;
  assign queue_bits_fu_op__T_4_en = io_enq_1_valid;
  assign queue_bits_fu_op__T_5_data = 5'h0;
  assign queue_bits_fu_op__T_5_addr = 6'h0;
  assign queue_bits_fu_op__T_5_mask = 1'h0;
  assign queue_bits_fu_op__T_5_en = 1'h0;
  assign queue_bits_fu_op__T_6_data = 5'h0;
  assign queue_bits_fu_op__T_6_addr = 6'h1;
  assign queue_bits_fu_op__T_6_mask = 1'h0;
  assign queue_bits_fu_op__T_6_en = 1'h0;
  assign queue_bits_fu_op__T_7_data = 5'h0;
  assign queue_bits_fu_op__T_7_addr = 6'h2;
  assign queue_bits_fu_op__T_7_mask = 1'h0;
  assign queue_bits_fu_op__T_7_en = 1'h0;
  assign queue_bits_fu_op__T_8_data = 5'h0;
  assign queue_bits_fu_op__T_8_addr = 6'h3;
  assign queue_bits_fu_op__T_8_mask = 1'h0;
  assign queue_bits_fu_op__T_8_en = 1'h0;
  assign queue_bits_fu_op__T_9_data = 5'h0;
  assign queue_bits_fu_op__T_9_addr = 6'h4;
  assign queue_bits_fu_op__T_9_mask = 1'h0;
  assign queue_bits_fu_op__T_9_en = 1'h0;
  assign queue_bits_fu_op__T_10_data = 5'h0;
  assign queue_bits_fu_op__T_10_addr = 6'h5;
  assign queue_bits_fu_op__T_10_mask = 1'h0;
  assign queue_bits_fu_op__T_10_en = 1'h0;
  assign queue_bits_fu_op__T_11_data = 5'h0;
  assign queue_bits_fu_op__T_11_addr = 6'h6;
  assign queue_bits_fu_op__T_11_mask = 1'h0;
  assign queue_bits_fu_op__T_11_en = 1'h0;
  assign queue_bits_fu_op__T_12_data = 5'h0;
  assign queue_bits_fu_op__T_12_addr = 6'h7;
  assign queue_bits_fu_op__T_12_mask = 1'h0;
  assign queue_bits_fu_op__T_12_en = 1'h0;
  assign queue_bits_fu_op__T_13_data = 5'h0;
  assign queue_bits_fu_op__T_13_addr = 6'h8;
  assign queue_bits_fu_op__T_13_mask = 1'h0;
  assign queue_bits_fu_op__T_13_en = 1'h0;
  assign queue_bits_fu_op__T_14_data = 5'h0;
  assign queue_bits_fu_op__T_14_addr = 6'h9;
  assign queue_bits_fu_op__T_14_mask = 1'h0;
  assign queue_bits_fu_op__T_14_en = 1'h0;
  assign queue_bits_fu_op__T_15_data = 5'h0;
  assign queue_bits_fu_op__T_15_addr = 6'ha;
  assign queue_bits_fu_op__T_15_mask = 1'h0;
  assign queue_bits_fu_op__T_15_en = 1'h0;
  assign queue_bits_fu_op__T_16_data = 5'h0;
  assign queue_bits_fu_op__T_16_addr = 6'hb;
  assign queue_bits_fu_op__T_16_mask = 1'h0;
  assign queue_bits_fu_op__T_16_en = 1'h0;
  assign queue_bits_fu_op__T_17_data = 5'h0;
  assign queue_bits_fu_op__T_17_addr = 6'hc;
  assign queue_bits_fu_op__T_17_mask = 1'h0;
  assign queue_bits_fu_op__T_17_en = 1'h0;
  assign queue_bits_fu_op__T_18_data = 5'h0;
  assign queue_bits_fu_op__T_18_addr = 6'hd;
  assign queue_bits_fu_op__T_18_mask = 1'h0;
  assign queue_bits_fu_op__T_18_en = 1'h0;
  assign queue_bits_fu_op__T_19_data = 5'h0;
  assign queue_bits_fu_op__T_19_addr = 6'he;
  assign queue_bits_fu_op__T_19_mask = 1'h0;
  assign queue_bits_fu_op__T_19_en = 1'h0;
  assign queue_bits_fu_op__T_20_data = 5'h0;
  assign queue_bits_fu_op__T_20_addr = 6'hf;
  assign queue_bits_fu_op__T_20_mask = 1'h0;
  assign queue_bits_fu_op__T_20_en = 1'h0;
  assign queue_bits_fu_op__T_21_data = 5'h0;
  assign queue_bits_fu_op__T_21_addr = 6'h10;
  assign queue_bits_fu_op__T_21_mask = 1'h0;
  assign queue_bits_fu_op__T_21_en = 1'h0;
  assign queue_bits_fu_op__T_22_data = 5'h0;
  assign queue_bits_fu_op__T_22_addr = 6'h11;
  assign queue_bits_fu_op__T_22_mask = 1'h0;
  assign queue_bits_fu_op__T_22_en = 1'h0;
  assign queue_bits_fu_op__T_23_data = 5'h0;
  assign queue_bits_fu_op__T_23_addr = 6'h12;
  assign queue_bits_fu_op__T_23_mask = 1'h0;
  assign queue_bits_fu_op__T_23_en = 1'h0;
  assign queue_bits_fu_op__T_24_data = 5'h0;
  assign queue_bits_fu_op__T_24_addr = 6'h13;
  assign queue_bits_fu_op__T_24_mask = 1'h0;
  assign queue_bits_fu_op__T_24_en = 1'h0;
  assign queue_bits_fu_op__T_25_data = 5'h0;
  assign queue_bits_fu_op__T_25_addr = 6'h14;
  assign queue_bits_fu_op__T_25_mask = 1'h0;
  assign queue_bits_fu_op__T_25_en = 1'h0;
  assign queue_bits_fu_op__T_26_data = 5'h0;
  assign queue_bits_fu_op__T_26_addr = 6'h15;
  assign queue_bits_fu_op__T_26_mask = 1'h0;
  assign queue_bits_fu_op__T_26_en = 1'h0;
  assign queue_bits_fu_op__T_27_data = 5'h0;
  assign queue_bits_fu_op__T_27_addr = 6'h16;
  assign queue_bits_fu_op__T_27_mask = 1'h0;
  assign queue_bits_fu_op__T_27_en = 1'h0;
  assign queue_bits_fu_op__T_28_data = 5'h0;
  assign queue_bits_fu_op__T_28_addr = 6'h17;
  assign queue_bits_fu_op__T_28_mask = 1'h0;
  assign queue_bits_fu_op__T_28_en = 1'h0;
  assign queue_bits_fu_op__T_29_data = 5'h0;
  assign queue_bits_fu_op__T_29_addr = 6'h18;
  assign queue_bits_fu_op__T_29_mask = 1'h0;
  assign queue_bits_fu_op__T_29_en = 1'h0;
  assign queue_bits_fu_op__T_30_data = 5'h0;
  assign queue_bits_fu_op__T_30_addr = 6'h19;
  assign queue_bits_fu_op__T_30_mask = 1'h0;
  assign queue_bits_fu_op__T_30_en = 1'h0;
  assign queue_bits_fu_op__T_31_data = 5'h0;
  assign queue_bits_fu_op__T_31_addr = 6'h1a;
  assign queue_bits_fu_op__T_31_mask = 1'h0;
  assign queue_bits_fu_op__T_31_en = 1'h0;
  assign queue_bits_fu_op__T_32_data = 5'h0;
  assign queue_bits_fu_op__T_32_addr = 6'h1b;
  assign queue_bits_fu_op__T_32_mask = 1'h0;
  assign queue_bits_fu_op__T_32_en = 1'h0;
  assign queue_bits_fu_op__T_33_data = 5'h0;
  assign queue_bits_fu_op__T_33_addr = 6'h1c;
  assign queue_bits_fu_op__T_33_mask = 1'h0;
  assign queue_bits_fu_op__T_33_en = 1'h0;
  assign queue_bits_fu_op__T_34_data = 5'h0;
  assign queue_bits_fu_op__T_34_addr = 6'h1d;
  assign queue_bits_fu_op__T_34_mask = 1'h0;
  assign queue_bits_fu_op__T_34_en = 1'h0;
  assign queue_bits_fu_op__T_35_data = 5'h0;
  assign queue_bits_fu_op__T_35_addr = 6'h1e;
  assign queue_bits_fu_op__T_35_mask = 1'h0;
  assign queue_bits_fu_op__T_35_en = 1'h0;
  assign queue_bits_fu_op__T_36_data = 5'h0;
  assign queue_bits_fu_op__T_36_addr = 6'h1f;
  assign queue_bits_fu_op__T_36_mask = 1'h0;
  assign queue_bits_fu_op__T_36_en = 1'h0;
  assign queue_bits_fu_op__T_37_data = 5'h0;
  assign queue_bits_fu_op__T_37_addr = 6'h20;
  assign queue_bits_fu_op__T_37_mask = 1'h0;
  assign queue_bits_fu_op__T_37_en = 1'h0;
  assign queue_bits_fu_op__T_38_data = 5'h0;
  assign queue_bits_fu_op__T_38_addr = 6'h21;
  assign queue_bits_fu_op__T_38_mask = 1'h0;
  assign queue_bits_fu_op__T_38_en = 1'h0;
  assign queue_bits_fu_op__T_39_data = 5'h0;
  assign queue_bits_fu_op__T_39_addr = 6'h22;
  assign queue_bits_fu_op__T_39_mask = 1'h0;
  assign queue_bits_fu_op__T_39_en = 1'h0;
  assign queue_bits_fu_op__T_40_data = 5'h0;
  assign queue_bits_fu_op__T_40_addr = 6'h23;
  assign queue_bits_fu_op__T_40_mask = 1'h0;
  assign queue_bits_fu_op__T_40_en = 1'h0;
  assign queue_bits_fu_op__T_41_data = 5'h0;
  assign queue_bits_fu_op__T_41_addr = 6'h24;
  assign queue_bits_fu_op__T_41_mask = 1'h0;
  assign queue_bits_fu_op__T_41_en = 1'h0;
  assign queue_bits_fu_op__T_42_data = 5'h0;
  assign queue_bits_fu_op__T_42_addr = 6'h25;
  assign queue_bits_fu_op__T_42_mask = 1'h0;
  assign queue_bits_fu_op__T_42_en = 1'h0;
  assign queue_bits_fu_op__T_43_data = 5'h0;
  assign queue_bits_fu_op__T_43_addr = 6'h26;
  assign queue_bits_fu_op__T_43_mask = 1'h0;
  assign queue_bits_fu_op__T_43_en = 1'h0;
  assign queue_bits_fu_op__T_44_data = 5'h0;
  assign queue_bits_fu_op__T_44_addr = 6'h27;
  assign queue_bits_fu_op__T_44_mask = 1'h0;
  assign queue_bits_fu_op__T_44_en = 1'h0;
  assign queue_bits_fu_op__T_45_data = 5'h0;
  assign queue_bits_fu_op__T_45_addr = 6'h28;
  assign queue_bits_fu_op__T_45_mask = 1'h0;
  assign queue_bits_fu_op__T_45_en = 1'h0;
  assign queue_bits_fu_op__T_46_data = 5'h0;
  assign queue_bits_fu_op__T_46_addr = 6'h29;
  assign queue_bits_fu_op__T_46_mask = 1'h0;
  assign queue_bits_fu_op__T_46_en = 1'h0;
  assign queue_bits_fu_op__T_47_data = 5'h0;
  assign queue_bits_fu_op__T_47_addr = 6'h2a;
  assign queue_bits_fu_op__T_47_mask = 1'h0;
  assign queue_bits_fu_op__T_47_en = 1'h0;
  assign queue_bits_fu_op__T_48_data = 5'h0;
  assign queue_bits_fu_op__T_48_addr = 6'h2b;
  assign queue_bits_fu_op__T_48_mask = 1'h0;
  assign queue_bits_fu_op__T_48_en = 1'h0;
  assign queue_bits_fu_op__T_49_data = 5'h0;
  assign queue_bits_fu_op__T_49_addr = 6'h2c;
  assign queue_bits_fu_op__T_49_mask = 1'h0;
  assign queue_bits_fu_op__T_49_en = 1'h0;
  assign queue_bits_fu_op__T_50_data = 5'h0;
  assign queue_bits_fu_op__T_50_addr = 6'h2d;
  assign queue_bits_fu_op__T_50_mask = 1'h0;
  assign queue_bits_fu_op__T_50_en = 1'h0;
  assign queue_bits_fu_op__T_51_data = 5'h0;
  assign queue_bits_fu_op__T_51_addr = 6'h2e;
  assign queue_bits_fu_op__T_51_mask = 1'h0;
  assign queue_bits_fu_op__T_51_en = 1'h0;
  assign queue_bits_fu_op__T_52_data = 5'h0;
  assign queue_bits_fu_op__T_52_addr = 6'h2f;
  assign queue_bits_fu_op__T_52_mask = 1'h0;
  assign queue_bits_fu_op__T_52_en = 1'h0;
  assign queue_bits_fu_op__T_53_data = 5'h0;
  assign queue_bits_fu_op__T_53_addr = 6'h30;
  assign queue_bits_fu_op__T_53_mask = 1'h0;
  assign queue_bits_fu_op__T_53_en = 1'h0;
  assign queue_bits_fu_op__T_54_data = 5'h0;
  assign queue_bits_fu_op__T_54_addr = 6'h31;
  assign queue_bits_fu_op__T_54_mask = 1'h0;
  assign queue_bits_fu_op__T_54_en = 1'h0;
  assign queue_bits_fu_op__T_55_data = 5'h0;
  assign queue_bits_fu_op__T_55_addr = 6'h32;
  assign queue_bits_fu_op__T_55_mask = 1'h0;
  assign queue_bits_fu_op__T_55_en = 1'h0;
  assign queue_bits_fu_op__T_56_data = 5'h0;
  assign queue_bits_fu_op__T_56_addr = 6'h33;
  assign queue_bits_fu_op__T_56_mask = 1'h0;
  assign queue_bits_fu_op__T_56_en = 1'h0;
  assign queue_bits_fu_op__T_57_data = 5'h0;
  assign queue_bits_fu_op__T_57_addr = 6'h34;
  assign queue_bits_fu_op__T_57_mask = 1'h0;
  assign queue_bits_fu_op__T_57_en = 1'h0;
  assign queue_bits_fu_op__T_58_data = 5'h0;
  assign queue_bits_fu_op__T_58_addr = 6'h35;
  assign queue_bits_fu_op__T_58_mask = 1'h0;
  assign queue_bits_fu_op__T_58_en = 1'h0;
  assign queue_bits_fu_op__T_59_data = 5'h0;
  assign queue_bits_fu_op__T_59_addr = 6'h36;
  assign queue_bits_fu_op__T_59_mask = 1'h0;
  assign queue_bits_fu_op__T_59_en = 1'h0;
  assign queue_bits_fu_op__T_60_data = 5'h0;
  assign queue_bits_fu_op__T_60_addr = 6'h37;
  assign queue_bits_fu_op__T_60_mask = 1'h0;
  assign queue_bits_fu_op__T_60_en = 1'h0;
  assign queue_bits_fu_op__T_61_data = 5'h0;
  assign queue_bits_fu_op__T_61_addr = 6'h38;
  assign queue_bits_fu_op__T_61_mask = 1'h0;
  assign queue_bits_fu_op__T_61_en = 1'h0;
  assign queue_bits_fu_op__T_62_data = 5'h0;
  assign queue_bits_fu_op__T_62_addr = 6'h39;
  assign queue_bits_fu_op__T_62_mask = 1'h0;
  assign queue_bits_fu_op__T_62_en = 1'h0;
  assign queue_bits_fu_op__T_63_data = 5'h0;
  assign queue_bits_fu_op__T_63_addr = 6'h3a;
  assign queue_bits_fu_op__T_63_mask = 1'h0;
  assign queue_bits_fu_op__T_63_en = 1'h0;
  assign queue_bits_fu_op__T_64_data = 5'h0;
  assign queue_bits_fu_op__T_64_addr = 6'h3b;
  assign queue_bits_fu_op__T_64_mask = 1'h0;
  assign queue_bits_fu_op__T_64_en = 1'h0;
  assign queue_bits_fu_op__T_65_data = 5'h0;
  assign queue_bits_fu_op__T_65_addr = 6'h3c;
  assign queue_bits_fu_op__T_65_mask = 1'h0;
  assign queue_bits_fu_op__T_65_en = 1'h0;
  assign queue_bits_fu_op__T_66_data = 5'h0;
  assign queue_bits_fu_op__T_66_addr = 6'h3d;
  assign queue_bits_fu_op__T_66_mask = 1'h0;
  assign queue_bits_fu_op__T_66_en = 1'h0;
  assign queue_bits_fu_op__T_67_data = 5'h0;
  assign queue_bits_fu_op__T_67_addr = 6'h3e;
  assign queue_bits_fu_op__T_67_mask = 1'h0;
  assign queue_bits_fu_op__T_67_en = 1'h0;
  assign queue_bits_fu_op__T_68_data = 5'h0;
  assign queue_bits_fu_op__T_68_addr = 6'h3f;
  assign queue_bits_fu_op__T_68_mask = 1'h0;
  assign queue_bits_fu_op__T_68_en = 1'h0;
  assign queue_bits_fu_op__T_70_data = 5'h0;
  assign queue_bits_fu_op__T_70_addr = 6'h0;
  assign queue_bits_fu_op__T_70_mask = 1'h0;
  assign queue_bits_fu_op__T_70_en = reset;
  assign queue_bits_fu_op__T_71_data = 5'h0;
  assign queue_bits_fu_op__T_71_addr = 6'h1;
  assign queue_bits_fu_op__T_71_mask = 1'h0;
  assign queue_bits_fu_op__T_71_en = reset;
  assign queue_bits_fu_op__T_72_data = 5'h0;
  assign queue_bits_fu_op__T_72_addr = 6'h2;
  assign queue_bits_fu_op__T_72_mask = 1'h0;
  assign queue_bits_fu_op__T_72_en = reset;
  assign queue_bits_fu_op__T_73_data = 5'h0;
  assign queue_bits_fu_op__T_73_addr = 6'h3;
  assign queue_bits_fu_op__T_73_mask = 1'h0;
  assign queue_bits_fu_op__T_73_en = reset;
  assign queue_bits_fu_op__T_74_data = 5'h0;
  assign queue_bits_fu_op__T_74_addr = 6'h4;
  assign queue_bits_fu_op__T_74_mask = 1'h0;
  assign queue_bits_fu_op__T_74_en = reset;
  assign queue_bits_fu_op__T_75_data = 5'h0;
  assign queue_bits_fu_op__T_75_addr = 6'h5;
  assign queue_bits_fu_op__T_75_mask = 1'h0;
  assign queue_bits_fu_op__T_75_en = reset;
  assign queue_bits_fu_op__T_76_data = 5'h0;
  assign queue_bits_fu_op__T_76_addr = 6'h6;
  assign queue_bits_fu_op__T_76_mask = 1'h0;
  assign queue_bits_fu_op__T_76_en = reset;
  assign queue_bits_fu_op__T_77_data = 5'h0;
  assign queue_bits_fu_op__T_77_addr = 6'h7;
  assign queue_bits_fu_op__T_77_mask = 1'h0;
  assign queue_bits_fu_op__T_77_en = reset;
  assign queue_bits_fu_op__T_78_data = 5'h0;
  assign queue_bits_fu_op__T_78_addr = 6'h8;
  assign queue_bits_fu_op__T_78_mask = 1'h0;
  assign queue_bits_fu_op__T_78_en = reset;
  assign queue_bits_fu_op__T_79_data = 5'h0;
  assign queue_bits_fu_op__T_79_addr = 6'h9;
  assign queue_bits_fu_op__T_79_mask = 1'h0;
  assign queue_bits_fu_op__T_79_en = reset;
  assign queue_bits_fu_op__T_80_data = 5'h0;
  assign queue_bits_fu_op__T_80_addr = 6'ha;
  assign queue_bits_fu_op__T_80_mask = 1'h0;
  assign queue_bits_fu_op__T_80_en = reset;
  assign queue_bits_fu_op__T_81_data = 5'h0;
  assign queue_bits_fu_op__T_81_addr = 6'hb;
  assign queue_bits_fu_op__T_81_mask = 1'h0;
  assign queue_bits_fu_op__T_81_en = reset;
  assign queue_bits_fu_op__T_82_data = 5'h0;
  assign queue_bits_fu_op__T_82_addr = 6'hc;
  assign queue_bits_fu_op__T_82_mask = 1'h0;
  assign queue_bits_fu_op__T_82_en = reset;
  assign queue_bits_fu_op__T_83_data = 5'h0;
  assign queue_bits_fu_op__T_83_addr = 6'hd;
  assign queue_bits_fu_op__T_83_mask = 1'h0;
  assign queue_bits_fu_op__T_83_en = reset;
  assign queue_bits_fu_op__T_84_data = 5'h0;
  assign queue_bits_fu_op__T_84_addr = 6'he;
  assign queue_bits_fu_op__T_84_mask = 1'h0;
  assign queue_bits_fu_op__T_84_en = reset;
  assign queue_bits_fu_op__T_85_data = 5'h0;
  assign queue_bits_fu_op__T_85_addr = 6'hf;
  assign queue_bits_fu_op__T_85_mask = 1'h0;
  assign queue_bits_fu_op__T_85_en = reset;
  assign queue_bits_fu_op__T_86_data = 5'h0;
  assign queue_bits_fu_op__T_86_addr = 6'h10;
  assign queue_bits_fu_op__T_86_mask = 1'h0;
  assign queue_bits_fu_op__T_86_en = reset;
  assign queue_bits_fu_op__T_87_data = 5'h0;
  assign queue_bits_fu_op__T_87_addr = 6'h11;
  assign queue_bits_fu_op__T_87_mask = 1'h0;
  assign queue_bits_fu_op__T_87_en = reset;
  assign queue_bits_fu_op__T_88_data = 5'h0;
  assign queue_bits_fu_op__T_88_addr = 6'h12;
  assign queue_bits_fu_op__T_88_mask = 1'h0;
  assign queue_bits_fu_op__T_88_en = reset;
  assign queue_bits_fu_op__T_89_data = 5'h0;
  assign queue_bits_fu_op__T_89_addr = 6'h13;
  assign queue_bits_fu_op__T_89_mask = 1'h0;
  assign queue_bits_fu_op__T_89_en = reset;
  assign queue_bits_fu_op__T_90_data = 5'h0;
  assign queue_bits_fu_op__T_90_addr = 6'h14;
  assign queue_bits_fu_op__T_90_mask = 1'h0;
  assign queue_bits_fu_op__T_90_en = reset;
  assign queue_bits_fu_op__T_91_data = 5'h0;
  assign queue_bits_fu_op__T_91_addr = 6'h15;
  assign queue_bits_fu_op__T_91_mask = 1'h0;
  assign queue_bits_fu_op__T_91_en = reset;
  assign queue_bits_fu_op__T_92_data = 5'h0;
  assign queue_bits_fu_op__T_92_addr = 6'h16;
  assign queue_bits_fu_op__T_92_mask = 1'h0;
  assign queue_bits_fu_op__T_92_en = reset;
  assign queue_bits_fu_op__T_93_data = 5'h0;
  assign queue_bits_fu_op__T_93_addr = 6'h17;
  assign queue_bits_fu_op__T_93_mask = 1'h0;
  assign queue_bits_fu_op__T_93_en = reset;
  assign queue_bits_fu_op__T_94_data = 5'h0;
  assign queue_bits_fu_op__T_94_addr = 6'h18;
  assign queue_bits_fu_op__T_94_mask = 1'h0;
  assign queue_bits_fu_op__T_94_en = reset;
  assign queue_bits_fu_op__T_95_data = 5'h0;
  assign queue_bits_fu_op__T_95_addr = 6'h19;
  assign queue_bits_fu_op__T_95_mask = 1'h0;
  assign queue_bits_fu_op__T_95_en = reset;
  assign queue_bits_fu_op__T_96_data = 5'h0;
  assign queue_bits_fu_op__T_96_addr = 6'h1a;
  assign queue_bits_fu_op__T_96_mask = 1'h0;
  assign queue_bits_fu_op__T_96_en = reset;
  assign queue_bits_fu_op__T_97_data = 5'h0;
  assign queue_bits_fu_op__T_97_addr = 6'h1b;
  assign queue_bits_fu_op__T_97_mask = 1'h0;
  assign queue_bits_fu_op__T_97_en = reset;
  assign queue_bits_fu_op__T_98_data = 5'h0;
  assign queue_bits_fu_op__T_98_addr = 6'h1c;
  assign queue_bits_fu_op__T_98_mask = 1'h0;
  assign queue_bits_fu_op__T_98_en = reset;
  assign queue_bits_fu_op__T_99_data = 5'h0;
  assign queue_bits_fu_op__T_99_addr = 6'h1d;
  assign queue_bits_fu_op__T_99_mask = 1'h0;
  assign queue_bits_fu_op__T_99_en = reset;
  assign queue_bits_fu_op__T_100_data = 5'h0;
  assign queue_bits_fu_op__T_100_addr = 6'h1e;
  assign queue_bits_fu_op__T_100_mask = 1'h0;
  assign queue_bits_fu_op__T_100_en = reset;
  assign queue_bits_fu_op__T_101_data = 5'h0;
  assign queue_bits_fu_op__T_101_addr = 6'h1f;
  assign queue_bits_fu_op__T_101_mask = 1'h0;
  assign queue_bits_fu_op__T_101_en = reset;
  assign queue_bits_fu_op__T_102_data = 5'h0;
  assign queue_bits_fu_op__T_102_addr = 6'h20;
  assign queue_bits_fu_op__T_102_mask = 1'h0;
  assign queue_bits_fu_op__T_102_en = reset;
  assign queue_bits_fu_op__T_103_data = 5'h0;
  assign queue_bits_fu_op__T_103_addr = 6'h21;
  assign queue_bits_fu_op__T_103_mask = 1'h0;
  assign queue_bits_fu_op__T_103_en = reset;
  assign queue_bits_fu_op__T_104_data = 5'h0;
  assign queue_bits_fu_op__T_104_addr = 6'h22;
  assign queue_bits_fu_op__T_104_mask = 1'h0;
  assign queue_bits_fu_op__T_104_en = reset;
  assign queue_bits_fu_op__T_105_data = 5'h0;
  assign queue_bits_fu_op__T_105_addr = 6'h23;
  assign queue_bits_fu_op__T_105_mask = 1'h0;
  assign queue_bits_fu_op__T_105_en = reset;
  assign queue_bits_fu_op__T_106_data = 5'h0;
  assign queue_bits_fu_op__T_106_addr = 6'h24;
  assign queue_bits_fu_op__T_106_mask = 1'h0;
  assign queue_bits_fu_op__T_106_en = reset;
  assign queue_bits_fu_op__T_107_data = 5'h0;
  assign queue_bits_fu_op__T_107_addr = 6'h25;
  assign queue_bits_fu_op__T_107_mask = 1'h0;
  assign queue_bits_fu_op__T_107_en = reset;
  assign queue_bits_fu_op__T_108_data = 5'h0;
  assign queue_bits_fu_op__T_108_addr = 6'h26;
  assign queue_bits_fu_op__T_108_mask = 1'h0;
  assign queue_bits_fu_op__T_108_en = reset;
  assign queue_bits_fu_op__T_109_data = 5'h0;
  assign queue_bits_fu_op__T_109_addr = 6'h27;
  assign queue_bits_fu_op__T_109_mask = 1'h0;
  assign queue_bits_fu_op__T_109_en = reset;
  assign queue_bits_fu_op__T_110_data = 5'h0;
  assign queue_bits_fu_op__T_110_addr = 6'h28;
  assign queue_bits_fu_op__T_110_mask = 1'h0;
  assign queue_bits_fu_op__T_110_en = reset;
  assign queue_bits_fu_op__T_111_data = 5'h0;
  assign queue_bits_fu_op__T_111_addr = 6'h29;
  assign queue_bits_fu_op__T_111_mask = 1'h0;
  assign queue_bits_fu_op__T_111_en = reset;
  assign queue_bits_fu_op__T_112_data = 5'h0;
  assign queue_bits_fu_op__T_112_addr = 6'h2a;
  assign queue_bits_fu_op__T_112_mask = 1'h0;
  assign queue_bits_fu_op__T_112_en = reset;
  assign queue_bits_fu_op__T_113_data = 5'h0;
  assign queue_bits_fu_op__T_113_addr = 6'h2b;
  assign queue_bits_fu_op__T_113_mask = 1'h0;
  assign queue_bits_fu_op__T_113_en = reset;
  assign queue_bits_fu_op__T_114_data = 5'h0;
  assign queue_bits_fu_op__T_114_addr = 6'h2c;
  assign queue_bits_fu_op__T_114_mask = 1'h0;
  assign queue_bits_fu_op__T_114_en = reset;
  assign queue_bits_fu_op__T_115_data = 5'h0;
  assign queue_bits_fu_op__T_115_addr = 6'h2d;
  assign queue_bits_fu_op__T_115_mask = 1'h0;
  assign queue_bits_fu_op__T_115_en = reset;
  assign queue_bits_fu_op__T_116_data = 5'h0;
  assign queue_bits_fu_op__T_116_addr = 6'h2e;
  assign queue_bits_fu_op__T_116_mask = 1'h0;
  assign queue_bits_fu_op__T_116_en = reset;
  assign queue_bits_fu_op__T_117_data = 5'h0;
  assign queue_bits_fu_op__T_117_addr = 6'h2f;
  assign queue_bits_fu_op__T_117_mask = 1'h0;
  assign queue_bits_fu_op__T_117_en = reset;
  assign queue_bits_fu_op__T_118_data = 5'h0;
  assign queue_bits_fu_op__T_118_addr = 6'h30;
  assign queue_bits_fu_op__T_118_mask = 1'h0;
  assign queue_bits_fu_op__T_118_en = reset;
  assign queue_bits_fu_op__T_119_data = 5'h0;
  assign queue_bits_fu_op__T_119_addr = 6'h31;
  assign queue_bits_fu_op__T_119_mask = 1'h0;
  assign queue_bits_fu_op__T_119_en = reset;
  assign queue_bits_fu_op__T_120_data = 5'h0;
  assign queue_bits_fu_op__T_120_addr = 6'h32;
  assign queue_bits_fu_op__T_120_mask = 1'h0;
  assign queue_bits_fu_op__T_120_en = reset;
  assign queue_bits_fu_op__T_121_data = 5'h0;
  assign queue_bits_fu_op__T_121_addr = 6'h33;
  assign queue_bits_fu_op__T_121_mask = 1'h0;
  assign queue_bits_fu_op__T_121_en = reset;
  assign queue_bits_fu_op__T_122_data = 5'h0;
  assign queue_bits_fu_op__T_122_addr = 6'h34;
  assign queue_bits_fu_op__T_122_mask = 1'h0;
  assign queue_bits_fu_op__T_122_en = reset;
  assign queue_bits_fu_op__T_123_data = 5'h0;
  assign queue_bits_fu_op__T_123_addr = 6'h35;
  assign queue_bits_fu_op__T_123_mask = 1'h0;
  assign queue_bits_fu_op__T_123_en = reset;
  assign queue_bits_fu_op__T_124_data = 5'h0;
  assign queue_bits_fu_op__T_124_addr = 6'h36;
  assign queue_bits_fu_op__T_124_mask = 1'h0;
  assign queue_bits_fu_op__T_124_en = reset;
  assign queue_bits_fu_op__T_125_data = 5'h0;
  assign queue_bits_fu_op__T_125_addr = 6'h37;
  assign queue_bits_fu_op__T_125_mask = 1'h0;
  assign queue_bits_fu_op__T_125_en = reset;
  assign queue_bits_fu_op__T_126_data = 5'h0;
  assign queue_bits_fu_op__T_126_addr = 6'h38;
  assign queue_bits_fu_op__T_126_mask = 1'h0;
  assign queue_bits_fu_op__T_126_en = reset;
  assign queue_bits_fu_op__T_127_data = 5'h0;
  assign queue_bits_fu_op__T_127_addr = 6'h39;
  assign queue_bits_fu_op__T_127_mask = 1'h0;
  assign queue_bits_fu_op__T_127_en = reset;
  assign queue_bits_fu_op__T_128_data = 5'h0;
  assign queue_bits_fu_op__T_128_addr = 6'h3a;
  assign queue_bits_fu_op__T_128_mask = 1'h0;
  assign queue_bits_fu_op__T_128_en = reset;
  assign queue_bits_fu_op__T_129_data = 5'h0;
  assign queue_bits_fu_op__T_129_addr = 6'h3b;
  assign queue_bits_fu_op__T_129_mask = 1'h0;
  assign queue_bits_fu_op__T_129_en = reset;
  assign queue_bits_fu_op__T_130_data = 5'h0;
  assign queue_bits_fu_op__T_130_addr = 6'h3c;
  assign queue_bits_fu_op__T_130_mask = 1'h0;
  assign queue_bits_fu_op__T_130_en = reset;
  assign queue_bits_fu_op__T_131_data = 5'h0;
  assign queue_bits_fu_op__T_131_addr = 6'h3d;
  assign queue_bits_fu_op__T_131_mask = 1'h0;
  assign queue_bits_fu_op__T_131_en = reset;
  assign queue_bits_fu_op__T_132_data = 5'h0;
  assign queue_bits_fu_op__T_132_addr = 6'h3e;
  assign queue_bits_fu_op__T_132_mask = 1'h0;
  assign queue_bits_fu_op__T_132_en = reset;
  assign queue_bits_fu_op__T_133_data = 5'h0;
  assign queue_bits_fu_op__T_133_addr = 6'h3f;
  assign queue_bits_fu_op__T_133_mask = 1'h0;
  assign queue_bits_fu_op__T_133_en = reset;
  assign queue_bits_fu_op_q_head_w_data = 5'h0;
  assign queue_bits_fu_op_q_head_w_addr = head;
  assign queue_bits_fu_op_q_head_w_mask = 1'h0;
  assign queue_bits_fu_op_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_id_q_head_r_addr = head;
  assign queue_bits_wb_id_q_head_r_data = queue_bits_wb_id[queue_bits_wb_id_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_id__T_3_data = io_enq_0_bits_data_wb_id;
  assign queue_bits_wb_id__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_id__T_3_mask = 1'h1;
  assign queue_bits_wb_id__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_id__T_4_data = io_enq_1_bits_data_wb_id;
  assign queue_bits_wb_id__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_id__T_4_mask = 1'h1;
  assign queue_bits_wb_id__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_id__T_5_data = 8'h0;
  assign queue_bits_wb_id__T_5_addr = 6'h0;
  assign queue_bits_wb_id__T_5_mask = 1'h0;
  assign queue_bits_wb_id__T_5_en = 1'h0;
  assign queue_bits_wb_id__T_6_data = 8'h0;
  assign queue_bits_wb_id__T_6_addr = 6'h1;
  assign queue_bits_wb_id__T_6_mask = 1'h0;
  assign queue_bits_wb_id__T_6_en = 1'h0;
  assign queue_bits_wb_id__T_7_data = 8'h0;
  assign queue_bits_wb_id__T_7_addr = 6'h2;
  assign queue_bits_wb_id__T_7_mask = 1'h0;
  assign queue_bits_wb_id__T_7_en = 1'h0;
  assign queue_bits_wb_id__T_8_data = 8'h0;
  assign queue_bits_wb_id__T_8_addr = 6'h3;
  assign queue_bits_wb_id__T_8_mask = 1'h0;
  assign queue_bits_wb_id__T_8_en = 1'h0;
  assign queue_bits_wb_id__T_9_data = 8'h0;
  assign queue_bits_wb_id__T_9_addr = 6'h4;
  assign queue_bits_wb_id__T_9_mask = 1'h0;
  assign queue_bits_wb_id__T_9_en = 1'h0;
  assign queue_bits_wb_id__T_10_data = 8'h0;
  assign queue_bits_wb_id__T_10_addr = 6'h5;
  assign queue_bits_wb_id__T_10_mask = 1'h0;
  assign queue_bits_wb_id__T_10_en = 1'h0;
  assign queue_bits_wb_id__T_11_data = 8'h0;
  assign queue_bits_wb_id__T_11_addr = 6'h6;
  assign queue_bits_wb_id__T_11_mask = 1'h0;
  assign queue_bits_wb_id__T_11_en = 1'h0;
  assign queue_bits_wb_id__T_12_data = 8'h0;
  assign queue_bits_wb_id__T_12_addr = 6'h7;
  assign queue_bits_wb_id__T_12_mask = 1'h0;
  assign queue_bits_wb_id__T_12_en = 1'h0;
  assign queue_bits_wb_id__T_13_data = 8'h0;
  assign queue_bits_wb_id__T_13_addr = 6'h8;
  assign queue_bits_wb_id__T_13_mask = 1'h0;
  assign queue_bits_wb_id__T_13_en = 1'h0;
  assign queue_bits_wb_id__T_14_data = 8'h0;
  assign queue_bits_wb_id__T_14_addr = 6'h9;
  assign queue_bits_wb_id__T_14_mask = 1'h0;
  assign queue_bits_wb_id__T_14_en = 1'h0;
  assign queue_bits_wb_id__T_15_data = 8'h0;
  assign queue_bits_wb_id__T_15_addr = 6'ha;
  assign queue_bits_wb_id__T_15_mask = 1'h0;
  assign queue_bits_wb_id__T_15_en = 1'h0;
  assign queue_bits_wb_id__T_16_data = 8'h0;
  assign queue_bits_wb_id__T_16_addr = 6'hb;
  assign queue_bits_wb_id__T_16_mask = 1'h0;
  assign queue_bits_wb_id__T_16_en = 1'h0;
  assign queue_bits_wb_id__T_17_data = 8'h0;
  assign queue_bits_wb_id__T_17_addr = 6'hc;
  assign queue_bits_wb_id__T_17_mask = 1'h0;
  assign queue_bits_wb_id__T_17_en = 1'h0;
  assign queue_bits_wb_id__T_18_data = 8'h0;
  assign queue_bits_wb_id__T_18_addr = 6'hd;
  assign queue_bits_wb_id__T_18_mask = 1'h0;
  assign queue_bits_wb_id__T_18_en = 1'h0;
  assign queue_bits_wb_id__T_19_data = 8'h0;
  assign queue_bits_wb_id__T_19_addr = 6'he;
  assign queue_bits_wb_id__T_19_mask = 1'h0;
  assign queue_bits_wb_id__T_19_en = 1'h0;
  assign queue_bits_wb_id__T_20_data = 8'h0;
  assign queue_bits_wb_id__T_20_addr = 6'hf;
  assign queue_bits_wb_id__T_20_mask = 1'h0;
  assign queue_bits_wb_id__T_20_en = 1'h0;
  assign queue_bits_wb_id__T_21_data = 8'h0;
  assign queue_bits_wb_id__T_21_addr = 6'h10;
  assign queue_bits_wb_id__T_21_mask = 1'h0;
  assign queue_bits_wb_id__T_21_en = 1'h0;
  assign queue_bits_wb_id__T_22_data = 8'h0;
  assign queue_bits_wb_id__T_22_addr = 6'h11;
  assign queue_bits_wb_id__T_22_mask = 1'h0;
  assign queue_bits_wb_id__T_22_en = 1'h0;
  assign queue_bits_wb_id__T_23_data = 8'h0;
  assign queue_bits_wb_id__T_23_addr = 6'h12;
  assign queue_bits_wb_id__T_23_mask = 1'h0;
  assign queue_bits_wb_id__T_23_en = 1'h0;
  assign queue_bits_wb_id__T_24_data = 8'h0;
  assign queue_bits_wb_id__T_24_addr = 6'h13;
  assign queue_bits_wb_id__T_24_mask = 1'h0;
  assign queue_bits_wb_id__T_24_en = 1'h0;
  assign queue_bits_wb_id__T_25_data = 8'h0;
  assign queue_bits_wb_id__T_25_addr = 6'h14;
  assign queue_bits_wb_id__T_25_mask = 1'h0;
  assign queue_bits_wb_id__T_25_en = 1'h0;
  assign queue_bits_wb_id__T_26_data = 8'h0;
  assign queue_bits_wb_id__T_26_addr = 6'h15;
  assign queue_bits_wb_id__T_26_mask = 1'h0;
  assign queue_bits_wb_id__T_26_en = 1'h0;
  assign queue_bits_wb_id__T_27_data = 8'h0;
  assign queue_bits_wb_id__T_27_addr = 6'h16;
  assign queue_bits_wb_id__T_27_mask = 1'h0;
  assign queue_bits_wb_id__T_27_en = 1'h0;
  assign queue_bits_wb_id__T_28_data = 8'h0;
  assign queue_bits_wb_id__T_28_addr = 6'h17;
  assign queue_bits_wb_id__T_28_mask = 1'h0;
  assign queue_bits_wb_id__T_28_en = 1'h0;
  assign queue_bits_wb_id__T_29_data = 8'h0;
  assign queue_bits_wb_id__T_29_addr = 6'h18;
  assign queue_bits_wb_id__T_29_mask = 1'h0;
  assign queue_bits_wb_id__T_29_en = 1'h0;
  assign queue_bits_wb_id__T_30_data = 8'h0;
  assign queue_bits_wb_id__T_30_addr = 6'h19;
  assign queue_bits_wb_id__T_30_mask = 1'h0;
  assign queue_bits_wb_id__T_30_en = 1'h0;
  assign queue_bits_wb_id__T_31_data = 8'h0;
  assign queue_bits_wb_id__T_31_addr = 6'h1a;
  assign queue_bits_wb_id__T_31_mask = 1'h0;
  assign queue_bits_wb_id__T_31_en = 1'h0;
  assign queue_bits_wb_id__T_32_data = 8'h0;
  assign queue_bits_wb_id__T_32_addr = 6'h1b;
  assign queue_bits_wb_id__T_32_mask = 1'h0;
  assign queue_bits_wb_id__T_32_en = 1'h0;
  assign queue_bits_wb_id__T_33_data = 8'h0;
  assign queue_bits_wb_id__T_33_addr = 6'h1c;
  assign queue_bits_wb_id__T_33_mask = 1'h0;
  assign queue_bits_wb_id__T_33_en = 1'h0;
  assign queue_bits_wb_id__T_34_data = 8'h0;
  assign queue_bits_wb_id__T_34_addr = 6'h1d;
  assign queue_bits_wb_id__T_34_mask = 1'h0;
  assign queue_bits_wb_id__T_34_en = 1'h0;
  assign queue_bits_wb_id__T_35_data = 8'h0;
  assign queue_bits_wb_id__T_35_addr = 6'h1e;
  assign queue_bits_wb_id__T_35_mask = 1'h0;
  assign queue_bits_wb_id__T_35_en = 1'h0;
  assign queue_bits_wb_id__T_36_data = 8'h0;
  assign queue_bits_wb_id__T_36_addr = 6'h1f;
  assign queue_bits_wb_id__T_36_mask = 1'h0;
  assign queue_bits_wb_id__T_36_en = 1'h0;
  assign queue_bits_wb_id__T_37_data = 8'h0;
  assign queue_bits_wb_id__T_37_addr = 6'h20;
  assign queue_bits_wb_id__T_37_mask = 1'h0;
  assign queue_bits_wb_id__T_37_en = 1'h0;
  assign queue_bits_wb_id__T_38_data = 8'h0;
  assign queue_bits_wb_id__T_38_addr = 6'h21;
  assign queue_bits_wb_id__T_38_mask = 1'h0;
  assign queue_bits_wb_id__T_38_en = 1'h0;
  assign queue_bits_wb_id__T_39_data = 8'h0;
  assign queue_bits_wb_id__T_39_addr = 6'h22;
  assign queue_bits_wb_id__T_39_mask = 1'h0;
  assign queue_bits_wb_id__T_39_en = 1'h0;
  assign queue_bits_wb_id__T_40_data = 8'h0;
  assign queue_bits_wb_id__T_40_addr = 6'h23;
  assign queue_bits_wb_id__T_40_mask = 1'h0;
  assign queue_bits_wb_id__T_40_en = 1'h0;
  assign queue_bits_wb_id__T_41_data = 8'h0;
  assign queue_bits_wb_id__T_41_addr = 6'h24;
  assign queue_bits_wb_id__T_41_mask = 1'h0;
  assign queue_bits_wb_id__T_41_en = 1'h0;
  assign queue_bits_wb_id__T_42_data = 8'h0;
  assign queue_bits_wb_id__T_42_addr = 6'h25;
  assign queue_bits_wb_id__T_42_mask = 1'h0;
  assign queue_bits_wb_id__T_42_en = 1'h0;
  assign queue_bits_wb_id__T_43_data = 8'h0;
  assign queue_bits_wb_id__T_43_addr = 6'h26;
  assign queue_bits_wb_id__T_43_mask = 1'h0;
  assign queue_bits_wb_id__T_43_en = 1'h0;
  assign queue_bits_wb_id__T_44_data = 8'h0;
  assign queue_bits_wb_id__T_44_addr = 6'h27;
  assign queue_bits_wb_id__T_44_mask = 1'h0;
  assign queue_bits_wb_id__T_44_en = 1'h0;
  assign queue_bits_wb_id__T_45_data = 8'h0;
  assign queue_bits_wb_id__T_45_addr = 6'h28;
  assign queue_bits_wb_id__T_45_mask = 1'h0;
  assign queue_bits_wb_id__T_45_en = 1'h0;
  assign queue_bits_wb_id__T_46_data = 8'h0;
  assign queue_bits_wb_id__T_46_addr = 6'h29;
  assign queue_bits_wb_id__T_46_mask = 1'h0;
  assign queue_bits_wb_id__T_46_en = 1'h0;
  assign queue_bits_wb_id__T_47_data = 8'h0;
  assign queue_bits_wb_id__T_47_addr = 6'h2a;
  assign queue_bits_wb_id__T_47_mask = 1'h0;
  assign queue_bits_wb_id__T_47_en = 1'h0;
  assign queue_bits_wb_id__T_48_data = 8'h0;
  assign queue_bits_wb_id__T_48_addr = 6'h2b;
  assign queue_bits_wb_id__T_48_mask = 1'h0;
  assign queue_bits_wb_id__T_48_en = 1'h0;
  assign queue_bits_wb_id__T_49_data = 8'h0;
  assign queue_bits_wb_id__T_49_addr = 6'h2c;
  assign queue_bits_wb_id__T_49_mask = 1'h0;
  assign queue_bits_wb_id__T_49_en = 1'h0;
  assign queue_bits_wb_id__T_50_data = 8'h0;
  assign queue_bits_wb_id__T_50_addr = 6'h2d;
  assign queue_bits_wb_id__T_50_mask = 1'h0;
  assign queue_bits_wb_id__T_50_en = 1'h0;
  assign queue_bits_wb_id__T_51_data = 8'h0;
  assign queue_bits_wb_id__T_51_addr = 6'h2e;
  assign queue_bits_wb_id__T_51_mask = 1'h0;
  assign queue_bits_wb_id__T_51_en = 1'h0;
  assign queue_bits_wb_id__T_52_data = 8'h0;
  assign queue_bits_wb_id__T_52_addr = 6'h2f;
  assign queue_bits_wb_id__T_52_mask = 1'h0;
  assign queue_bits_wb_id__T_52_en = 1'h0;
  assign queue_bits_wb_id__T_53_data = 8'h0;
  assign queue_bits_wb_id__T_53_addr = 6'h30;
  assign queue_bits_wb_id__T_53_mask = 1'h0;
  assign queue_bits_wb_id__T_53_en = 1'h0;
  assign queue_bits_wb_id__T_54_data = 8'h0;
  assign queue_bits_wb_id__T_54_addr = 6'h31;
  assign queue_bits_wb_id__T_54_mask = 1'h0;
  assign queue_bits_wb_id__T_54_en = 1'h0;
  assign queue_bits_wb_id__T_55_data = 8'h0;
  assign queue_bits_wb_id__T_55_addr = 6'h32;
  assign queue_bits_wb_id__T_55_mask = 1'h0;
  assign queue_bits_wb_id__T_55_en = 1'h0;
  assign queue_bits_wb_id__T_56_data = 8'h0;
  assign queue_bits_wb_id__T_56_addr = 6'h33;
  assign queue_bits_wb_id__T_56_mask = 1'h0;
  assign queue_bits_wb_id__T_56_en = 1'h0;
  assign queue_bits_wb_id__T_57_data = 8'h0;
  assign queue_bits_wb_id__T_57_addr = 6'h34;
  assign queue_bits_wb_id__T_57_mask = 1'h0;
  assign queue_bits_wb_id__T_57_en = 1'h0;
  assign queue_bits_wb_id__T_58_data = 8'h0;
  assign queue_bits_wb_id__T_58_addr = 6'h35;
  assign queue_bits_wb_id__T_58_mask = 1'h0;
  assign queue_bits_wb_id__T_58_en = 1'h0;
  assign queue_bits_wb_id__T_59_data = 8'h0;
  assign queue_bits_wb_id__T_59_addr = 6'h36;
  assign queue_bits_wb_id__T_59_mask = 1'h0;
  assign queue_bits_wb_id__T_59_en = 1'h0;
  assign queue_bits_wb_id__T_60_data = 8'h0;
  assign queue_bits_wb_id__T_60_addr = 6'h37;
  assign queue_bits_wb_id__T_60_mask = 1'h0;
  assign queue_bits_wb_id__T_60_en = 1'h0;
  assign queue_bits_wb_id__T_61_data = 8'h0;
  assign queue_bits_wb_id__T_61_addr = 6'h38;
  assign queue_bits_wb_id__T_61_mask = 1'h0;
  assign queue_bits_wb_id__T_61_en = 1'h0;
  assign queue_bits_wb_id__T_62_data = 8'h0;
  assign queue_bits_wb_id__T_62_addr = 6'h39;
  assign queue_bits_wb_id__T_62_mask = 1'h0;
  assign queue_bits_wb_id__T_62_en = 1'h0;
  assign queue_bits_wb_id__T_63_data = 8'h0;
  assign queue_bits_wb_id__T_63_addr = 6'h3a;
  assign queue_bits_wb_id__T_63_mask = 1'h0;
  assign queue_bits_wb_id__T_63_en = 1'h0;
  assign queue_bits_wb_id__T_64_data = 8'h0;
  assign queue_bits_wb_id__T_64_addr = 6'h3b;
  assign queue_bits_wb_id__T_64_mask = 1'h0;
  assign queue_bits_wb_id__T_64_en = 1'h0;
  assign queue_bits_wb_id__T_65_data = 8'h0;
  assign queue_bits_wb_id__T_65_addr = 6'h3c;
  assign queue_bits_wb_id__T_65_mask = 1'h0;
  assign queue_bits_wb_id__T_65_en = 1'h0;
  assign queue_bits_wb_id__T_66_data = 8'h0;
  assign queue_bits_wb_id__T_66_addr = 6'h3d;
  assign queue_bits_wb_id__T_66_mask = 1'h0;
  assign queue_bits_wb_id__T_66_en = 1'h0;
  assign queue_bits_wb_id__T_67_data = 8'h0;
  assign queue_bits_wb_id__T_67_addr = 6'h3e;
  assign queue_bits_wb_id__T_67_mask = 1'h0;
  assign queue_bits_wb_id__T_67_en = 1'h0;
  assign queue_bits_wb_id__T_68_data = 8'h0;
  assign queue_bits_wb_id__T_68_addr = 6'h3f;
  assign queue_bits_wb_id__T_68_mask = 1'h0;
  assign queue_bits_wb_id__T_68_en = 1'h0;
  assign queue_bits_wb_id__T_70_data = 8'h0;
  assign queue_bits_wb_id__T_70_addr = 6'h0;
  assign queue_bits_wb_id__T_70_mask = 1'h0;
  assign queue_bits_wb_id__T_70_en = reset;
  assign queue_bits_wb_id__T_71_data = 8'h0;
  assign queue_bits_wb_id__T_71_addr = 6'h1;
  assign queue_bits_wb_id__T_71_mask = 1'h0;
  assign queue_bits_wb_id__T_71_en = reset;
  assign queue_bits_wb_id__T_72_data = 8'h0;
  assign queue_bits_wb_id__T_72_addr = 6'h2;
  assign queue_bits_wb_id__T_72_mask = 1'h0;
  assign queue_bits_wb_id__T_72_en = reset;
  assign queue_bits_wb_id__T_73_data = 8'h0;
  assign queue_bits_wb_id__T_73_addr = 6'h3;
  assign queue_bits_wb_id__T_73_mask = 1'h0;
  assign queue_bits_wb_id__T_73_en = reset;
  assign queue_bits_wb_id__T_74_data = 8'h0;
  assign queue_bits_wb_id__T_74_addr = 6'h4;
  assign queue_bits_wb_id__T_74_mask = 1'h0;
  assign queue_bits_wb_id__T_74_en = reset;
  assign queue_bits_wb_id__T_75_data = 8'h0;
  assign queue_bits_wb_id__T_75_addr = 6'h5;
  assign queue_bits_wb_id__T_75_mask = 1'h0;
  assign queue_bits_wb_id__T_75_en = reset;
  assign queue_bits_wb_id__T_76_data = 8'h0;
  assign queue_bits_wb_id__T_76_addr = 6'h6;
  assign queue_bits_wb_id__T_76_mask = 1'h0;
  assign queue_bits_wb_id__T_76_en = reset;
  assign queue_bits_wb_id__T_77_data = 8'h0;
  assign queue_bits_wb_id__T_77_addr = 6'h7;
  assign queue_bits_wb_id__T_77_mask = 1'h0;
  assign queue_bits_wb_id__T_77_en = reset;
  assign queue_bits_wb_id__T_78_data = 8'h0;
  assign queue_bits_wb_id__T_78_addr = 6'h8;
  assign queue_bits_wb_id__T_78_mask = 1'h0;
  assign queue_bits_wb_id__T_78_en = reset;
  assign queue_bits_wb_id__T_79_data = 8'h0;
  assign queue_bits_wb_id__T_79_addr = 6'h9;
  assign queue_bits_wb_id__T_79_mask = 1'h0;
  assign queue_bits_wb_id__T_79_en = reset;
  assign queue_bits_wb_id__T_80_data = 8'h0;
  assign queue_bits_wb_id__T_80_addr = 6'ha;
  assign queue_bits_wb_id__T_80_mask = 1'h0;
  assign queue_bits_wb_id__T_80_en = reset;
  assign queue_bits_wb_id__T_81_data = 8'h0;
  assign queue_bits_wb_id__T_81_addr = 6'hb;
  assign queue_bits_wb_id__T_81_mask = 1'h0;
  assign queue_bits_wb_id__T_81_en = reset;
  assign queue_bits_wb_id__T_82_data = 8'h0;
  assign queue_bits_wb_id__T_82_addr = 6'hc;
  assign queue_bits_wb_id__T_82_mask = 1'h0;
  assign queue_bits_wb_id__T_82_en = reset;
  assign queue_bits_wb_id__T_83_data = 8'h0;
  assign queue_bits_wb_id__T_83_addr = 6'hd;
  assign queue_bits_wb_id__T_83_mask = 1'h0;
  assign queue_bits_wb_id__T_83_en = reset;
  assign queue_bits_wb_id__T_84_data = 8'h0;
  assign queue_bits_wb_id__T_84_addr = 6'he;
  assign queue_bits_wb_id__T_84_mask = 1'h0;
  assign queue_bits_wb_id__T_84_en = reset;
  assign queue_bits_wb_id__T_85_data = 8'h0;
  assign queue_bits_wb_id__T_85_addr = 6'hf;
  assign queue_bits_wb_id__T_85_mask = 1'h0;
  assign queue_bits_wb_id__T_85_en = reset;
  assign queue_bits_wb_id__T_86_data = 8'h0;
  assign queue_bits_wb_id__T_86_addr = 6'h10;
  assign queue_bits_wb_id__T_86_mask = 1'h0;
  assign queue_bits_wb_id__T_86_en = reset;
  assign queue_bits_wb_id__T_87_data = 8'h0;
  assign queue_bits_wb_id__T_87_addr = 6'h11;
  assign queue_bits_wb_id__T_87_mask = 1'h0;
  assign queue_bits_wb_id__T_87_en = reset;
  assign queue_bits_wb_id__T_88_data = 8'h0;
  assign queue_bits_wb_id__T_88_addr = 6'h12;
  assign queue_bits_wb_id__T_88_mask = 1'h0;
  assign queue_bits_wb_id__T_88_en = reset;
  assign queue_bits_wb_id__T_89_data = 8'h0;
  assign queue_bits_wb_id__T_89_addr = 6'h13;
  assign queue_bits_wb_id__T_89_mask = 1'h0;
  assign queue_bits_wb_id__T_89_en = reset;
  assign queue_bits_wb_id__T_90_data = 8'h0;
  assign queue_bits_wb_id__T_90_addr = 6'h14;
  assign queue_bits_wb_id__T_90_mask = 1'h0;
  assign queue_bits_wb_id__T_90_en = reset;
  assign queue_bits_wb_id__T_91_data = 8'h0;
  assign queue_bits_wb_id__T_91_addr = 6'h15;
  assign queue_bits_wb_id__T_91_mask = 1'h0;
  assign queue_bits_wb_id__T_91_en = reset;
  assign queue_bits_wb_id__T_92_data = 8'h0;
  assign queue_bits_wb_id__T_92_addr = 6'h16;
  assign queue_bits_wb_id__T_92_mask = 1'h0;
  assign queue_bits_wb_id__T_92_en = reset;
  assign queue_bits_wb_id__T_93_data = 8'h0;
  assign queue_bits_wb_id__T_93_addr = 6'h17;
  assign queue_bits_wb_id__T_93_mask = 1'h0;
  assign queue_bits_wb_id__T_93_en = reset;
  assign queue_bits_wb_id__T_94_data = 8'h0;
  assign queue_bits_wb_id__T_94_addr = 6'h18;
  assign queue_bits_wb_id__T_94_mask = 1'h0;
  assign queue_bits_wb_id__T_94_en = reset;
  assign queue_bits_wb_id__T_95_data = 8'h0;
  assign queue_bits_wb_id__T_95_addr = 6'h19;
  assign queue_bits_wb_id__T_95_mask = 1'h0;
  assign queue_bits_wb_id__T_95_en = reset;
  assign queue_bits_wb_id__T_96_data = 8'h0;
  assign queue_bits_wb_id__T_96_addr = 6'h1a;
  assign queue_bits_wb_id__T_96_mask = 1'h0;
  assign queue_bits_wb_id__T_96_en = reset;
  assign queue_bits_wb_id__T_97_data = 8'h0;
  assign queue_bits_wb_id__T_97_addr = 6'h1b;
  assign queue_bits_wb_id__T_97_mask = 1'h0;
  assign queue_bits_wb_id__T_97_en = reset;
  assign queue_bits_wb_id__T_98_data = 8'h0;
  assign queue_bits_wb_id__T_98_addr = 6'h1c;
  assign queue_bits_wb_id__T_98_mask = 1'h0;
  assign queue_bits_wb_id__T_98_en = reset;
  assign queue_bits_wb_id__T_99_data = 8'h0;
  assign queue_bits_wb_id__T_99_addr = 6'h1d;
  assign queue_bits_wb_id__T_99_mask = 1'h0;
  assign queue_bits_wb_id__T_99_en = reset;
  assign queue_bits_wb_id__T_100_data = 8'h0;
  assign queue_bits_wb_id__T_100_addr = 6'h1e;
  assign queue_bits_wb_id__T_100_mask = 1'h0;
  assign queue_bits_wb_id__T_100_en = reset;
  assign queue_bits_wb_id__T_101_data = 8'h0;
  assign queue_bits_wb_id__T_101_addr = 6'h1f;
  assign queue_bits_wb_id__T_101_mask = 1'h0;
  assign queue_bits_wb_id__T_101_en = reset;
  assign queue_bits_wb_id__T_102_data = 8'h0;
  assign queue_bits_wb_id__T_102_addr = 6'h20;
  assign queue_bits_wb_id__T_102_mask = 1'h0;
  assign queue_bits_wb_id__T_102_en = reset;
  assign queue_bits_wb_id__T_103_data = 8'h0;
  assign queue_bits_wb_id__T_103_addr = 6'h21;
  assign queue_bits_wb_id__T_103_mask = 1'h0;
  assign queue_bits_wb_id__T_103_en = reset;
  assign queue_bits_wb_id__T_104_data = 8'h0;
  assign queue_bits_wb_id__T_104_addr = 6'h22;
  assign queue_bits_wb_id__T_104_mask = 1'h0;
  assign queue_bits_wb_id__T_104_en = reset;
  assign queue_bits_wb_id__T_105_data = 8'h0;
  assign queue_bits_wb_id__T_105_addr = 6'h23;
  assign queue_bits_wb_id__T_105_mask = 1'h0;
  assign queue_bits_wb_id__T_105_en = reset;
  assign queue_bits_wb_id__T_106_data = 8'h0;
  assign queue_bits_wb_id__T_106_addr = 6'h24;
  assign queue_bits_wb_id__T_106_mask = 1'h0;
  assign queue_bits_wb_id__T_106_en = reset;
  assign queue_bits_wb_id__T_107_data = 8'h0;
  assign queue_bits_wb_id__T_107_addr = 6'h25;
  assign queue_bits_wb_id__T_107_mask = 1'h0;
  assign queue_bits_wb_id__T_107_en = reset;
  assign queue_bits_wb_id__T_108_data = 8'h0;
  assign queue_bits_wb_id__T_108_addr = 6'h26;
  assign queue_bits_wb_id__T_108_mask = 1'h0;
  assign queue_bits_wb_id__T_108_en = reset;
  assign queue_bits_wb_id__T_109_data = 8'h0;
  assign queue_bits_wb_id__T_109_addr = 6'h27;
  assign queue_bits_wb_id__T_109_mask = 1'h0;
  assign queue_bits_wb_id__T_109_en = reset;
  assign queue_bits_wb_id__T_110_data = 8'h0;
  assign queue_bits_wb_id__T_110_addr = 6'h28;
  assign queue_bits_wb_id__T_110_mask = 1'h0;
  assign queue_bits_wb_id__T_110_en = reset;
  assign queue_bits_wb_id__T_111_data = 8'h0;
  assign queue_bits_wb_id__T_111_addr = 6'h29;
  assign queue_bits_wb_id__T_111_mask = 1'h0;
  assign queue_bits_wb_id__T_111_en = reset;
  assign queue_bits_wb_id__T_112_data = 8'h0;
  assign queue_bits_wb_id__T_112_addr = 6'h2a;
  assign queue_bits_wb_id__T_112_mask = 1'h0;
  assign queue_bits_wb_id__T_112_en = reset;
  assign queue_bits_wb_id__T_113_data = 8'h0;
  assign queue_bits_wb_id__T_113_addr = 6'h2b;
  assign queue_bits_wb_id__T_113_mask = 1'h0;
  assign queue_bits_wb_id__T_113_en = reset;
  assign queue_bits_wb_id__T_114_data = 8'h0;
  assign queue_bits_wb_id__T_114_addr = 6'h2c;
  assign queue_bits_wb_id__T_114_mask = 1'h0;
  assign queue_bits_wb_id__T_114_en = reset;
  assign queue_bits_wb_id__T_115_data = 8'h0;
  assign queue_bits_wb_id__T_115_addr = 6'h2d;
  assign queue_bits_wb_id__T_115_mask = 1'h0;
  assign queue_bits_wb_id__T_115_en = reset;
  assign queue_bits_wb_id__T_116_data = 8'h0;
  assign queue_bits_wb_id__T_116_addr = 6'h2e;
  assign queue_bits_wb_id__T_116_mask = 1'h0;
  assign queue_bits_wb_id__T_116_en = reset;
  assign queue_bits_wb_id__T_117_data = 8'h0;
  assign queue_bits_wb_id__T_117_addr = 6'h2f;
  assign queue_bits_wb_id__T_117_mask = 1'h0;
  assign queue_bits_wb_id__T_117_en = reset;
  assign queue_bits_wb_id__T_118_data = 8'h0;
  assign queue_bits_wb_id__T_118_addr = 6'h30;
  assign queue_bits_wb_id__T_118_mask = 1'h0;
  assign queue_bits_wb_id__T_118_en = reset;
  assign queue_bits_wb_id__T_119_data = 8'h0;
  assign queue_bits_wb_id__T_119_addr = 6'h31;
  assign queue_bits_wb_id__T_119_mask = 1'h0;
  assign queue_bits_wb_id__T_119_en = reset;
  assign queue_bits_wb_id__T_120_data = 8'h0;
  assign queue_bits_wb_id__T_120_addr = 6'h32;
  assign queue_bits_wb_id__T_120_mask = 1'h0;
  assign queue_bits_wb_id__T_120_en = reset;
  assign queue_bits_wb_id__T_121_data = 8'h0;
  assign queue_bits_wb_id__T_121_addr = 6'h33;
  assign queue_bits_wb_id__T_121_mask = 1'h0;
  assign queue_bits_wb_id__T_121_en = reset;
  assign queue_bits_wb_id__T_122_data = 8'h0;
  assign queue_bits_wb_id__T_122_addr = 6'h34;
  assign queue_bits_wb_id__T_122_mask = 1'h0;
  assign queue_bits_wb_id__T_122_en = reset;
  assign queue_bits_wb_id__T_123_data = 8'h0;
  assign queue_bits_wb_id__T_123_addr = 6'h35;
  assign queue_bits_wb_id__T_123_mask = 1'h0;
  assign queue_bits_wb_id__T_123_en = reset;
  assign queue_bits_wb_id__T_124_data = 8'h0;
  assign queue_bits_wb_id__T_124_addr = 6'h36;
  assign queue_bits_wb_id__T_124_mask = 1'h0;
  assign queue_bits_wb_id__T_124_en = reset;
  assign queue_bits_wb_id__T_125_data = 8'h0;
  assign queue_bits_wb_id__T_125_addr = 6'h37;
  assign queue_bits_wb_id__T_125_mask = 1'h0;
  assign queue_bits_wb_id__T_125_en = reset;
  assign queue_bits_wb_id__T_126_data = 8'h0;
  assign queue_bits_wb_id__T_126_addr = 6'h38;
  assign queue_bits_wb_id__T_126_mask = 1'h0;
  assign queue_bits_wb_id__T_126_en = reset;
  assign queue_bits_wb_id__T_127_data = 8'h0;
  assign queue_bits_wb_id__T_127_addr = 6'h39;
  assign queue_bits_wb_id__T_127_mask = 1'h0;
  assign queue_bits_wb_id__T_127_en = reset;
  assign queue_bits_wb_id__T_128_data = 8'h0;
  assign queue_bits_wb_id__T_128_addr = 6'h3a;
  assign queue_bits_wb_id__T_128_mask = 1'h0;
  assign queue_bits_wb_id__T_128_en = reset;
  assign queue_bits_wb_id__T_129_data = 8'h0;
  assign queue_bits_wb_id__T_129_addr = 6'h3b;
  assign queue_bits_wb_id__T_129_mask = 1'h0;
  assign queue_bits_wb_id__T_129_en = reset;
  assign queue_bits_wb_id__T_130_data = 8'h0;
  assign queue_bits_wb_id__T_130_addr = 6'h3c;
  assign queue_bits_wb_id__T_130_mask = 1'h0;
  assign queue_bits_wb_id__T_130_en = reset;
  assign queue_bits_wb_id__T_131_data = 8'h0;
  assign queue_bits_wb_id__T_131_addr = 6'h3d;
  assign queue_bits_wb_id__T_131_mask = 1'h0;
  assign queue_bits_wb_id__T_131_en = reset;
  assign queue_bits_wb_id__T_132_data = 8'h0;
  assign queue_bits_wb_id__T_132_addr = 6'h3e;
  assign queue_bits_wb_id__T_132_mask = 1'h0;
  assign queue_bits_wb_id__T_132_en = reset;
  assign queue_bits_wb_id__T_133_data = 8'h0;
  assign queue_bits_wb_id__T_133_addr = 6'h3f;
  assign queue_bits_wb_id__T_133_mask = 1'h0;
  assign queue_bits_wb_id__T_133_en = reset;
  assign queue_bits_wb_id_q_head_w_data = 8'h0;
  assign queue_bits_wb_id_q_head_w_addr = head;
  assign queue_bits_wb_id_q_head_w_mask = 1'h0;
  assign queue_bits_wb_id_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_pc_q_head_r_addr = head;
  assign queue_bits_wb_pc_q_head_r_data = queue_bits_wb_pc[queue_bits_wb_pc_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_pc__T_3_data = io_enq_0_bits_data_wb_pc;
  assign queue_bits_wb_pc__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_pc__T_3_mask = 1'h1;
  assign queue_bits_wb_pc__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_pc__T_4_data = io_enq_1_bits_data_wb_pc;
  assign queue_bits_wb_pc__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_pc__T_4_mask = 1'h1;
  assign queue_bits_wb_pc__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_pc__T_5_data = 32'h0;
  assign queue_bits_wb_pc__T_5_addr = 6'h0;
  assign queue_bits_wb_pc__T_5_mask = 1'h0;
  assign queue_bits_wb_pc__T_5_en = 1'h0;
  assign queue_bits_wb_pc__T_6_data = 32'h0;
  assign queue_bits_wb_pc__T_6_addr = 6'h1;
  assign queue_bits_wb_pc__T_6_mask = 1'h0;
  assign queue_bits_wb_pc__T_6_en = 1'h0;
  assign queue_bits_wb_pc__T_7_data = 32'h0;
  assign queue_bits_wb_pc__T_7_addr = 6'h2;
  assign queue_bits_wb_pc__T_7_mask = 1'h0;
  assign queue_bits_wb_pc__T_7_en = 1'h0;
  assign queue_bits_wb_pc__T_8_data = 32'h0;
  assign queue_bits_wb_pc__T_8_addr = 6'h3;
  assign queue_bits_wb_pc__T_8_mask = 1'h0;
  assign queue_bits_wb_pc__T_8_en = 1'h0;
  assign queue_bits_wb_pc__T_9_data = 32'h0;
  assign queue_bits_wb_pc__T_9_addr = 6'h4;
  assign queue_bits_wb_pc__T_9_mask = 1'h0;
  assign queue_bits_wb_pc__T_9_en = 1'h0;
  assign queue_bits_wb_pc__T_10_data = 32'h0;
  assign queue_bits_wb_pc__T_10_addr = 6'h5;
  assign queue_bits_wb_pc__T_10_mask = 1'h0;
  assign queue_bits_wb_pc__T_10_en = 1'h0;
  assign queue_bits_wb_pc__T_11_data = 32'h0;
  assign queue_bits_wb_pc__T_11_addr = 6'h6;
  assign queue_bits_wb_pc__T_11_mask = 1'h0;
  assign queue_bits_wb_pc__T_11_en = 1'h0;
  assign queue_bits_wb_pc__T_12_data = 32'h0;
  assign queue_bits_wb_pc__T_12_addr = 6'h7;
  assign queue_bits_wb_pc__T_12_mask = 1'h0;
  assign queue_bits_wb_pc__T_12_en = 1'h0;
  assign queue_bits_wb_pc__T_13_data = 32'h0;
  assign queue_bits_wb_pc__T_13_addr = 6'h8;
  assign queue_bits_wb_pc__T_13_mask = 1'h0;
  assign queue_bits_wb_pc__T_13_en = 1'h0;
  assign queue_bits_wb_pc__T_14_data = 32'h0;
  assign queue_bits_wb_pc__T_14_addr = 6'h9;
  assign queue_bits_wb_pc__T_14_mask = 1'h0;
  assign queue_bits_wb_pc__T_14_en = 1'h0;
  assign queue_bits_wb_pc__T_15_data = 32'h0;
  assign queue_bits_wb_pc__T_15_addr = 6'ha;
  assign queue_bits_wb_pc__T_15_mask = 1'h0;
  assign queue_bits_wb_pc__T_15_en = 1'h0;
  assign queue_bits_wb_pc__T_16_data = 32'h0;
  assign queue_bits_wb_pc__T_16_addr = 6'hb;
  assign queue_bits_wb_pc__T_16_mask = 1'h0;
  assign queue_bits_wb_pc__T_16_en = 1'h0;
  assign queue_bits_wb_pc__T_17_data = 32'h0;
  assign queue_bits_wb_pc__T_17_addr = 6'hc;
  assign queue_bits_wb_pc__T_17_mask = 1'h0;
  assign queue_bits_wb_pc__T_17_en = 1'h0;
  assign queue_bits_wb_pc__T_18_data = 32'h0;
  assign queue_bits_wb_pc__T_18_addr = 6'hd;
  assign queue_bits_wb_pc__T_18_mask = 1'h0;
  assign queue_bits_wb_pc__T_18_en = 1'h0;
  assign queue_bits_wb_pc__T_19_data = 32'h0;
  assign queue_bits_wb_pc__T_19_addr = 6'he;
  assign queue_bits_wb_pc__T_19_mask = 1'h0;
  assign queue_bits_wb_pc__T_19_en = 1'h0;
  assign queue_bits_wb_pc__T_20_data = 32'h0;
  assign queue_bits_wb_pc__T_20_addr = 6'hf;
  assign queue_bits_wb_pc__T_20_mask = 1'h0;
  assign queue_bits_wb_pc__T_20_en = 1'h0;
  assign queue_bits_wb_pc__T_21_data = 32'h0;
  assign queue_bits_wb_pc__T_21_addr = 6'h10;
  assign queue_bits_wb_pc__T_21_mask = 1'h0;
  assign queue_bits_wb_pc__T_21_en = 1'h0;
  assign queue_bits_wb_pc__T_22_data = 32'h0;
  assign queue_bits_wb_pc__T_22_addr = 6'h11;
  assign queue_bits_wb_pc__T_22_mask = 1'h0;
  assign queue_bits_wb_pc__T_22_en = 1'h0;
  assign queue_bits_wb_pc__T_23_data = 32'h0;
  assign queue_bits_wb_pc__T_23_addr = 6'h12;
  assign queue_bits_wb_pc__T_23_mask = 1'h0;
  assign queue_bits_wb_pc__T_23_en = 1'h0;
  assign queue_bits_wb_pc__T_24_data = 32'h0;
  assign queue_bits_wb_pc__T_24_addr = 6'h13;
  assign queue_bits_wb_pc__T_24_mask = 1'h0;
  assign queue_bits_wb_pc__T_24_en = 1'h0;
  assign queue_bits_wb_pc__T_25_data = 32'h0;
  assign queue_bits_wb_pc__T_25_addr = 6'h14;
  assign queue_bits_wb_pc__T_25_mask = 1'h0;
  assign queue_bits_wb_pc__T_25_en = 1'h0;
  assign queue_bits_wb_pc__T_26_data = 32'h0;
  assign queue_bits_wb_pc__T_26_addr = 6'h15;
  assign queue_bits_wb_pc__T_26_mask = 1'h0;
  assign queue_bits_wb_pc__T_26_en = 1'h0;
  assign queue_bits_wb_pc__T_27_data = 32'h0;
  assign queue_bits_wb_pc__T_27_addr = 6'h16;
  assign queue_bits_wb_pc__T_27_mask = 1'h0;
  assign queue_bits_wb_pc__T_27_en = 1'h0;
  assign queue_bits_wb_pc__T_28_data = 32'h0;
  assign queue_bits_wb_pc__T_28_addr = 6'h17;
  assign queue_bits_wb_pc__T_28_mask = 1'h0;
  assign queue_bits_wb_pc__T_28_en = 1'h0;
  assign queue_bits_wb_pc__T_29_data = 32'h0;
  assign queue_bits_wb_pc__T_29_addr = 6'h18;
  assign queue_bits_wb_pc__T_29_mask = 1'h0;
  assign queue_bits_wb_pc__T_29_en = 1'h0;
  assign queue_bits_wb_pc__T_30_data = 32'h0;
  assign queue_bits_wb_pc__T_30_addr = 6'h19;
  assign queue_bits_wb_pc__T_30_mask = 1'h0;
  assign queue_bits_wb_pc__T_30_en = 1'h0;
  assign queue_bits_wb_pc__T_31_data = 32'h0;
  assign queue_bits_wb_pc__T_31_addr = 6'h1a;
  assign queue_bits_wb_pc__T_31_mask = 1'h0;
  assign queue_bits_wb_pc__T_31_en = 1'h0;
  assign queue_bits_wb_pc__T_32_data = 32'h0;
  assign queue_bits_wb_pc__T_32_addr = 6'h1b;
  assign queue_bits_wb_pc__T_32_mask = 1'h0;
  assign queue_bits_wb_pc__T_32_en = 1'h0;
  assign queue_bits_wb_pc__T_33_data = 32'h0;
  assign queue_bits_wb_pc__T_33_addr = 6'h1c;
  assign queue_bits_wb_pc__T_33_mask = 1'h0;
  assign queue_bits_wb_pc__T_33_en = 1'h0;
  assign queue_bits_wb_pc__T_34_data = 32'h0;
  assign queue_bits_wb_pc__T_34_addr = 6'h1d;
  assign queue_bits_wb_pc__T_34_mask = 1'h0;
  assign queue_bits_wb_pc__T_34_en = 1'h0;
  assign queue_bits_wb_pc__T_35_data = 32'h0;
  assign queue_bits_wb_pc__T_35_addr = 6'h1e;
  assign queue_bits_wb_pc__T_35_mask = 1'h0;
  assign queue_bits_wb_pc__T_35_en = 1'h0;
  assign queue_bits_wb_pc__T_36_data = 32'h0;
  assign queue_bits_wb_pc__T_36_addr = 6'h1f;
  assign queue_bits_wb_pc__T_36_mask = 1'h0;
  assign queue_bits_wb_pc__T_36_en = 1'h0;
  assign queue_bits_wb_pc__T_37_data = 32'h0;
  assign queue_bits_wb_pc__T_37_addr = 6'h20;
  assign queue_bits_wb_pc__T_37_mask = 1'h0;
  assign queue_bits_wb_pc__T_37_en = 1'h0;
  assign queue_bits_wb_pc__T_38_data = 32'h0;
  assign queue_bits_wb_pc__T_38_addr = 6'h21;
  assign queue_bits_wb_pc__T_38_mask = 1'h0;
  assign queue_bits_wb_pc__T_38_en = 1'h0;
  assign queue_bits_wb_pc__T_39_data = 32'h0;
  assign queue_bits_wb_pc__T_39_addr = 6'h22;
  assign queue_bits_wb_pc__T_39_mask = 1'h0;
  assign queue_bits_wb_pc__T_39_en = 1'h0;
  assign queue_bits_wb_pc__T_40_data = 32'h0;
  assign queue_bits_wb_pc__T_40_addr = 6'h23;
  assign queue_bits_wb_pc__T_40_mask = 1'h0;
  assign queue_bits_wb_pc__T_40_en = 1'h0;
  assign queue_bits_wb_pc__T_41_data = 32'h0;
  assign queue_bits_wb_pc__T_41_addr = 6'h24;
  assign queue_bits_wb_pc__T_41_mask = 1'h0;
  assign queue_bits_wb_pc__T_41_en = 1'h0;
  assign queue_bits_wb_pc__T_42_data = 32'h0;
  assign queue_bits_wb_pc__T_42_addr = 6'h25;
  assign queue_bits_wb_pc__T_42_mask = 1'h0;
  assign queue_bits_wb_pc__T_42_en = 1'h0;
  assign queue_bits_wb_pc__T_43_data = 32'h0;
  assign queue_bits_wb_pc__T_43_addr = 6'h26;
  assign queue_bits_wb_pc__T_43_mask = 1'h0;
  assign queue_bits_wb_pc__T_43_en = 1'h0;
  assign queue_bits_wb_pc__T_44_data = 32'h0;
  assign queue_bits_wb_pc__T_44_addr = 6'h27;
  assign queue_bits_wb_pc__T_44_mask = 1'h0;
  assign queue_bits_wb_pc__T_44_en = 1'h0;
  assign queue_bits_wb_pc__T_45_data = 32'h0;
  assign queue_bits_wb_pc__T_45_addr = 6'h28;
  assign queue_bits_wb_pc__T_45_mask = 1'h0;
  assign queue_bits_wb_pc__T_45_en = 1'h0;
  assign queue_bits_wb_pc__T_46_data = 32'h0;
  assign queue_bits_wb_pc__T_46_addr = 6'h29;
  assign queue_bits_wb_pc__T_46_mask = 1'h0;
  assign queue_bits_wb_pc__T_46_en = 1'h0;
  assign queue_bits_wb_pc__T_47_data = 32'h0;
  assign queue_bits_wb_pc__T_47_addr = 6'h2a;
  assign queue_bits_wb_pc__T_47_mask = 1'h0;
  assign queue_bits_wb_pc__T_47_en = 1'h0;
  assign queue_bits_wb_pc__T_48_data = 32'h0;
  assign queue_bits_wb_pc__T_48_addr = 6'h2b;
  assign queue_bits_wb_pc__T_48_mask = 1'h0;
  assign queue_bits_wb_pc__T_48_en = 1'h0;
  assign queue_bits_wb_pc__T_49_data = 32'h0;
  assign queue_bits_wb_pc__T_49_addr = 6'h2c;
  assign queue_bits_wb_pc__T_49_mask = 1'h0;
  assign queue_bits_wb_pc__T_49_en = 1'h0;
  assign queue_bits_wb_pc__T_50_data = 32'h0;
  assign queue_bits_wb_pc__T_50_addr = 6'h2d;
  assign queue_bits_wb_pc__T_50_mask = 1'h0;
  assign queue_bits_wb_pc__T_50_en = 1'h0;
  assign queue_bits_wb_pc__T_51_data = 32'h0;
  assign queue_bits_wb_pc__T_51_addr = 6'h2e;
  assign queue_bits_wb_pc__T_51_mask = 1'h0;
  assign queue_bits_wb_pc__T_51_en = 1'h0;
  assign queue_bits_wb_pc__T_52_data = 32'h0;
  assign queue_bits_wb_pc__T_52_addr = 6'h2f;
  assign queue_bits_wb_pc__T_52_mask = 1'h0;
  assign queue_bits_wb_pc__T_52_en = 1'h0;
  assign queue_bits_wb_pc__T_53_data = 32'h0;
  assign queue_bits_wb_pc__T_53_addr = 6'h30;
  assign queue_bits_wb_pc__T_53_mask = 1'h0;
  assign queue_bits_wb_pc__T_53_en = 1'h0;
  assign queue_bits_wb_pc__T_54_data = 32'h0;
  assign queue_bits_wb_pc__T_54_addr = 6'h31;
  assign queue_bits_wb_pc__T_54_mask = 1'h0;
  assign queue_bits_wb_pc__T_54_en = 1'h0;
  assign queue_bits_wb_pc__T_55_data = 32'h0;
  assign queue_bits_wb_pc__T_55_addr = 6'h32;
  assign queue_bits_wb_pc__T_55_mask = 1'h0;
  assign queue_bits_wb_pc__T_55_en = 1'h0;
  assign queue_bits_wb_pc__T_56_data = 32'h0;
  assign queue_bits_wb_pc__T_56_addr = 6'h33;
  assign queue_bits_wb_pc__T_56_mask = 1'h0;
  assign queue_bits_wb_pc__T_56_en = 1'h0;
  assign queue_bits_wb_pc__T_57_data = 32'h0;
  assign queue_bits_wb_pc__T_57_addr = 6'h34;
  assign queue_bits_wb_pc__T_57_mask = 1'h0;
  assign queue_bits_wb_pc__T_57_en = 1'h0;
  assign queue_bits_wb_pc__T_58_data = 32'h0;
  assign queue_bits_wb_pc__T_58_addr = 6'h35;
  assign queue_bits_wb_pc__T_58_mask = 1'h0;
  assign queue_bits_wb_pc__T_58_en = 1'h0;
  assign queue_bits_wb_pc__T_59_data = 32'h0;
  assign queue_bits_wb_pc__T_59_addr = 6'h36;
  assign queue_bits_wb_pc__T_59_mask = 1'h0;
  assign queue_bits_wb_pc__T_59_en = 1'h0;
  assign queue_bits_wb_pc__T_60_data = 32'h0;
  assign queue_bits_wb_pc__T_60_addr = 6'h37;
  assign queue_bits_wb_pc__T_60_mask = 1'h0;
  assign queue_bits_wb_pc__T_60_en = 1'h0;
  assign queue_bits_wb_pc__T_61_data = 32'h0;
  assign queue_bits_wb_pc__T_61_addr = 6'h38;
  assign queue_bits_wb_pc__T_61_mask = 1'h0;
  assign queue_bits_wb_pc__T_61_en = 1'h0;
  assign queue_bits_wb_pc__T_62_data = 32'h0;
  assign queue_bits_wb_pc__T_62_addr = 6'h39;
  assign queue_bits_wb_pc__T_62_mask = 1'h0;
  assign queue_bits_wb_pc__T_62_en = 1'h0;
  assign queue_bits_wb_pc__T_63_data = 32'h0;
  assign queue_bits_wb_pc__T_63_addr = 6'h3a;
  assign queue_bits_wb_pc__T_63_mask = 1'h0;
  assign queue_bits_wb_pc__T_63_en = 1'h0;
  assign queue_bits_wb_pc__T_64_data = 32'h0;
  assign queue_bits_wb_pc__T_64_addr = 6'h3b;
  assign queue_bits_wb_pc__T_64_mask = 1'h0;
  assign queue_bits_wb_pc__T_64_en = 1'h0;
  assign queue_bits_wb_pc__T_65_data = 32'h0;
  assign queue_bits_wb_pc__T_65_addr = 6'h3c;
  assign queue_bits_wb_pc__T_65_mask = 1'h0;
  assign queue_bits_wb_pc__T_65_en = 1'h0;
  assign queue_bits_wb_pc__T_66_data = 32'h0;
  assign queue_bits_wb_pc__T_66_addr = 6'h3d;
  assign queue_bits_wb_pc__T_66_mask = 1'h0;
  assign queue_bits_wb_pc__T_66_en = 1'h0;
  assign queue_bits_wb_pc__T_67_data = 32'h0;
  assign queue_bits_wb_pc__T_67_addr = 6'h3e;
  assign queue_bits_wb_pc__T_67_mask = 1'h0;
  assign queue_bits_wb_pc__T_67_en = 1'h0;
  assign queue_bits_wb_pc__T_68_data = 32'h0;
  assign queue_bits_wb_pc__T_68_addr = 6'h3f;
  assign queue_bits_wb_pc__T_68_mask = 1'h0;
  assign queue_bits_wb_pc__T_68_en = 1'h0;
  assign queue_bits_wb_pc__T_70_data = 32'h0;
  assign queue_bits_wb_pc__T_70_addr = 6'h0;
  assign queue_bits_wb_pc__T_70_mask = 1'h0;
  assign queue_bits_wb_pc__T_70_en = reset;
  assign queue_bits_wb_pc__T_71_data = 32'h0;
  assign queue_bits_wb_pc__T_71_addr = 6'h1;
  assign queue_bits_wb_pc__T_71_mask = 1'h0;
  assign queue_bits_wb_pc__T_71_en = reset;
  assign queue_bits_wb_pc__T_72_data = 32'h0;
  assign queue_bits_wb_pc__T_72_addr = 6'h2;
  assign queue_bits_wb_pc__T_72_mask = 1'h0;
  assign queue_bits_wb_pc__T_72_en = reset;
  assign queue_bits_wb_pc__T_73_data = 32'h0;
  assign queue_bits_wb_pc__T_73_addr = 6'h3;
  assign queue_bits_wb_pc__T_73_mask = 1'h0;
  assign queue_bits_wb_pc__T_73_en = reset;
  assign queue_bits_wb_pc__T_74_data = 32'h0;
  assign queue_bits_wb_pc__T_74_addr = 6'h4;
  assign queue_bits_wb_pc__T_74_mask = 1'h0;
  assign queue_bits_wb_pc__T_74_en = reset;
  assign queue_bits_wb_pc__T_75_data = 32'h0;
  assign queue_bits_wb_pc__T_75_addr = 6'h5;
  assign queue_bits_wb_pc__T_75_mask = 1'h0;
  assign queue_bits_wb_pc__T_75_en = reset;
  assign queue_bits_wb_pc__T_76_data = 32'h0;
  assign queue_bits_wb_pc__T_76_addr = 6'h6;
  assign queue_bits_wb_pc__T_76_mask = 1'h0;
  assign queue_bits_wb_pc__T_76_en = reset;
  assign queue_bits_wb_pc__T_77_data = 32'h0;
  assign queue_bits_wb_pc__T_77_addr = 6'h7;
  assign queue_bits_wb_pc__T_77_mask = 1'h0;
  assign queue_bits_wb_pc__T_77_en = reset;
  assign queue_bits_wb_pc__T_78_data = 32'h0;
  assign queue_bits_wb_pc__T_78_addr = 6'h8;
  assign queue_bits_wb_pc__T_78_mask = 1'h0;
  assign queue_bits_wb_pc__T_78_en = reset;
  assign queue_bits_wb_pc__T_79_data = 32'h0;
  assign queue_bits_wb_pc__T_79_addr = 6'h9;
  assign queue_bits_wb_pc__T_79_mask = 1'h0;
  assign queue_bits_wb_pc__T_79_en = reset;
  assign queue_bits_wb_pc__T_80_data = 32'h0;
  assign queue_bits_wb_pc__T_80_addr = 6'ha;
  assign queue_bits_wb_pc__T_80_mask = 1'h0;
  assign queue_bits_wb_pc__T_80_en = reset;
  assign queue_bits_wb_pc__T_81_data = 32'h0;
  assign queue_bits_wb_pc__T_81_addr = 6'hb;
  assign queue_bits_wb_pc__T_81_mask = 1'h0;
  assign queue_bits_wb_pc__T_81_en = reset;
  assign queue_bits_wb_pc__T_82_data = 32'h0;
  assign queue_bits_wb_pc__T_82_addr = 6'hc;
  assign queue_bits_wb_pc__T_82_mask = 1'h0;
  assign queue_bits_wb_pc__T_82_en = reset;
  assign queue_bits_wb_pc__T_83_data = 32'h0;
  assign queue_bits_wb_pc__T_83_addr = 6'hd;
  assign queue_bits_wb_pc__T_83_mask = 1'h0;
  assign queue_bits_wb_pc__T_83_en = reset;
  assign queue_bits_wb_pc__T_84_data = 32'h0;
  assign queue_bits_wb_pc__T_84_addr = 6'he;
  assign queue_bits_wb_pc__T_84_mask = 1'h0;
  assign queue_bits_wb_pc__T_84_en = reset;
  assign queue_bits_wb_pc__T_85_data = 32'h0;
  assign queue_bits_wb_pc__T_85_addr = 6'hf;
  assign queue_bits_wb_pc__T_85_mask = 1'h0;
  assign queue_bits_wb_pc__T_85_en = reset;
  assign queue_bits_wb_pc__T_86_data = 32'h0;
  assign queue_bits_wb_pc__T_86_addr = 6'h10;
  assign queue_bits_wb_pc__T_86_mask = 1'h0;
  assign queue_bits_wb_pc__T_86_en = reset;
  assign queue_bits_wb_pc__T_87_data = 32'h0;
  assign queue_bits_wb_pc__T_87_addr = 6'h11;
  assign queue_bits_wb_pc__T_87_mask = 1'h0;
  assign queue_bits_wb_pc__T_87_en = reset;
  assign queue_bits_wb_pc__T_88_data = 32'h0;
  assign queue_bits_wb_pc__T_88_addr = 6'h12;
  assign queue_bits_wb_pc__T_88_mask = 1'h0;
  assign queue_bits_wb_pc__T_88_en = reset;
  assign queue_bits_wb_pc__T_89_data = 32'h0;
  assign queue_bits_wb_pc__T_89_addr = 6'h13;
  assign queue_bits_wb_pc__T_89_mask = 1'h0;
  assign queue_bits_wb_pc__T_89_en = reset;
  assign queue_bits_wb_pc__T_90_data = 32'h0;
  assign queue_bits_wb_pc__T_90_addr = 6'h14;
  assign queue_bits_wb_pc__T_90_mask = 1'h0;
  assign queue_bits_wb_pc__T_90_en = reset;
  assign queue_bits_wb_pc__T_91_data = 32'h0;
  assign queue_bits_wb_pc__T_91_addr = 6'h15;
  assign queue_bits_wb_pc__T_91_mask = 1'h0;
  assign queue_bits_wb_pc__T_91_en = reset;
  assign queue_bits_wb_pc__T_92_data = 32'h0;
  assign queue_bits_wb_pc__T_92_addr = 6'h16;
  assign queue_bits_wb_pc__T_92_mask = 1'h0;
  assign queue_bits_wb_pc__T_92_en = reset;
  assign queue_bits_wb_pc__T_93_data = 32'h0;
  assign queue_bits_wb_pc__T_93_addr = 6'h17;
  assign queue_bits_wb_pc__T_93_mask = 1'h0;
  assign queue_bits_wb_pc__T_93_en = reset;
  assign queue_bits_wb_pc__T_94_data = 32'h0;
  assign queue_bits_wb_pc__T_94_addr = 6'h18;
  assign queue_bits_wb_pc__T_94_mask = 1'h0;
  assign queue_bits_wb_pc__T_94_en = reset;
  assign queue_bits_wb_pc__T_95_data = 32'h0;
  assign queue_bits_wb_pc__T_95_addr = 6'h19;
  assign queue_bits_wb_pc__T_95_mask = 1'h0;
  assign queue_bits_wb_pc__T_95_en = reset;
  assign queue_bits_wb_pc__T_96_data = 32'h0;
  assign queue_bits_wb_pc__T_96_addr = 6'h1a;
  assign queue_bits_wb_pc__T_96_mask = 1'h0;
  assign queue_bits_wb_pc__T_96_en = reset;
  assign queue_bits_wb_pc__T_97_data = 32'h0;
  assign queue_bits_wb_pc__T_97_addr = 6'h1b;
  assign queue_bits_wb_pc__T_97_mask = 1'h0;
  assign queue_bits_wb_pc__T_97_en = reset;
  assign queue_bits_wb_pc__T_98_data = 32'h0;
  assign queue_bits_wb_pc__T_98_addr = 6'h1c;
  assign queue_bits_wb_pc__T_98_mask = 1'h0;
  assign queue_bits_wb_pc__T_98_en = reset;
  assign queue_bits_wb_pc__T_99_data = 32'h0;
  assign queue_bits_wb_pc__T_99_addr = 6'h1d;
  assign queue_bits_wb_pc__T_99_mask = 1'h0;
  assign queue_bits_wb_pc__T_99_en = reset;
  assign queue_bits_wb_pc__T_100_data = 32'h0;
  assign queue_bits_wb_pc__T_100_addr = 6'h1e;
  assign queue_bits_wb_pc__T_100_mask = 1'h0;
  assign queue_bits_wb_pc__T_100_en = reset;
  assign queue_bits_wb_pc__T_101_data = 32'h0;
  assign queue_bits_wb_pc__T_101_addr = 6'h1f;
  assign queue_bits_wb_pc__T_101_mask = 1'h0;
  assign queue_bits_wb_pc__T_101_en = reset;
  assign queue_bits_wb_pc__T_102_data = 32'h0;
  assign queue_bits_wb_pc__T_102_addr = 6'h20;
  assign queue_bits_wb_pc__T_102_mask = 1'h0;
  assign queue_bits_wb_pc__T_102_en = reset;
  assign queue_bits_wb_pc__T_103_data = 32'h0;
  assign queue_bits_wb_pc__T_103_addr = 6'h21;
  assign queue_bits_wb_pc__T_103_mask = 1'h0;
  assign queue_bits_wb_pc__T_103_en = reset;
  assign queue_bits_wb_pc__T_104_data = 32'h0;
  assign queue_bits_wb_pc__T_104_addr = 6'h22;
  assign queue_bits_wb_pc__T_104_mask = 1'h0;
  assign queue_bits_wb_pc__T_104_en = reset;
  assign queue_bits_wb_pc__T_105_data = 32'h0;
  assign queue_bits_wb_pc__T_105_addr = 6'h23;
  assign queue_bits_wb_pc__T_105_mask = 1'h0;
  assign queue_bits_wb_pc__T_105_en = reset;
  assign queue_bits_wb_pc__T_106_data = 32'h0;
  assign queue_bits_wb_pc__T_106_addr = 6'h24;
  assign queue_bits_wb_pc__T_106_mask = 1'h0;
  assign queue_bits_wb_pc__T_106_en = reset;
  assign queue_bits_wb_pc__T_107_data = 32'h0;
  assign queue_bits_wb_pc__T_107_addr = 6'h25;
  assign queue_bits_wb_pc__T_107_mask = 1'h0;
  assign queue_bits_wb_pc__T_107_en = reset;
  assign queue_bits_wb_pc__T_108_data = 32'h0;
  assign queue_bits_wb_pc__T_108_addr = 6'h26;
  assign queue_bits_wb_pc__T_108_mask = 1'h0;
  assign queue_bits_wb_pc__T_108_en = reset;
  assign queue_bits_wb_pc__T_109_data = 32'h0;
  assign queue_bits_wb_pc__T_109_addr = 6'h27;
  assign queue_bits_wb_pc__T_109_mask = 1'h0;
  assign queue_bits_wb_pc__T_109_en = reset;
  assign queue_bits_wb_pc__T_110_data = 32'h0;
  assign queue_bits_wb_pc__T_110_addr = 6'h28;
  assign queue_bits_wb_pc__T_110_mask = 1'h0;
  assign queue_bits_wb_pc__T_110_en = reset;
  assign queue_bits_wb_pc__T_111_data = 32'h0;
  assign queue_bits_wb_pc__T_111_addr = 6'h29;
  assign queue_bits_wb_pc__T_111_mask = 1'h0;
  assign queue_bits_wb_pc__T_111_en = reset;
  assign queue_bits_wb_pc__T_112_data = 32'h0;
  assign queue_bits_wb_pc__T_112_addr = 6'h2a;
  assign queue_bits_wb_pc__T_112_mask = 1'h0;
  assign queue_bits_wb_pc__T_112_en = reset;
  assign queue_bits_wb_pc__T_113_data = 32'h0;
  assign queue_bits_wb_pc__T_113_addr = 6'h2b;
  assign queue_bits_wb_pc__T_113_mask = 1'h0;
  assign queue_bits_wb_pc__T_113_en = reset;
  assign queue_bits_wb_pc__T_114_data = 32'h0;
  assign queue_bits_wb_pc__T_114_addr = 6'h2c;
  assign queue_bits_wb_pc__T_114_mask = 1'h0;
  assign queue_bits_wb_pc__T_114_en = reset;
  assign queue_bits_wb_pc__T_115_data = 32'h0;
  assign queue_bits_wb_pc__T_115_addr = 6'h2d;
  assign queue_bits_wb_pc__T_115_mask = 1'h0;
  assign queue_bits_wb_pc__T_115_en = reset;
  assign queue_bits_wb_pc__T_116_data = 32'h0;
  assign queue_bits_wb_pc__T_116_addr = 6'h2e;
  assign queue_bits_wb_pc__T_116_mask = 1'h0;
  assign queue_bits_wb_pc__T_116_en = reset;
  assign queue_bits_wb_pc__T_117_data = 32'h0;
  assign queue_bits_wb_pc__T_117_addr = 6'h2f;
  assign queue_bits_wb_pc__T_117_mask = 1'h0;
  assign queue_bits_wb_pc__T_117_en = reset;
  assign queue_bits_wb_pc__T_118_data = 32'h0;
  assign queue_bits_wb_pc__T_118_addr = 6'h30;
  assign queue_bits_wb_pc__T_118_mask = 1'h0;
  assign queue_bits_wb_pc__T_118_en = reset;
  assign queue_bits_wb_pc__T_119_data = 32'h0;
  assign queue_bits_wb_pc__T_119_addr = 6'h31;
  assign queue_bits_wb_pc__T_119_mask = 1'h0;
  assign queue_bits_wb_pc__T_119_en = reset;
  assign queue_bits_wb_pc__T_120_data = 32'h0;
  assign queue_bits_wb_pc__T_120_addr = 6'h32;
  assign queue_bits_wb_pc__T_120_mask = 1'h0;
  assign queue_bits_wb_pc__T_120_en = reset;
  assign queue_bits_wb_pc__T_121_data = 32'h0;
  assign queue_bits_wb_pc__T_121_addr = 6'h33;
  assign queue_bits_wb_pc__T_121_mask = 1'h0;
  assign queue_bits_wb_pc__T_121_en = reset;
  assign queue_bits_wb_pc__T_122_data = 32'h0;
  assign queue_bits_wb_pc__T_122_addr = 6'h34;
  assign queue_bits_wb_pc__T_122_mask = 1'h0;
  assign queue_bits_wb_pc__T_122_en = reset;
  assign queue_bits_wb_pc__T_123_data = 32'h0;
  assign queue_bits_wb_pc__T_123_addr = 6'h35;
  assign queue_bits_wb_pc__T_123_mask = 1'h0;
  assign queue_bits_wb_pc__T_123_en = reset;
  assign queue_bits_wb_pc__T_124_data = 32'h0;
  assign queue_bits_wb_pc__T_124_addr = 6'h36;
  assign queue_bits_wb_pc__T_124_mask = 1'h0;
  assign queue_bits_wb_pc__T_124_en = reset;
  assign queue_bits_wb_pc__T_125_data = 32'h0;
  assign queue_bits_wb_pc__T_125_addr = 6'h37;
  assign queue_bits_wb_pc__T_125_mask = 1'h0;
  assign queue_bits_wb_pc__T_125_en = reset;
  assign queue_bits_wb_pc__T_126_data = 32'h0;
  assign queue_bits_wb_pc__T_126_addr = 6'h38;
  assign queue_bits_wb_pc__T_126_mask = 1'h0;
  assign queue_bits_wb_pc__T_126_en = reset;
  assign queue_bits_wb_pc__T_127_data = 32'h0;
  assign queue_bits_wb_pc__T_127_addr = 6'h39;
  assign queue_bits_wb_pc__T_127_mask = 1'h0;
  assign queue_bits_wb_pc__T_127_en = reset;
  assign queue_bits_wb_pc__T_128_data = 32'h0;
  assign queue_bits_wb_pc__T_128_addr = 6'h3a;
  assign queue_bits_wb_pc__T_128_mask = 1'h0;
  assign queue_bits_wb_pc__T_128_en = reset;
  assign queue_bits_wb_pc__T_129_data = 32'h0;
  assign queue_bits_wb_pc__T_129_addr = 6'h3b;
  assign queue_bits_wb_pc__T_129_mask = 1'h0;
  assign queue_bits_wb_pc__T_129_en = reset;
  assign queue_bits_wb_pc__T_130_data = 32'h0;
  assign queue_bits_wb_pc__T_130_addr = 6'h3c;
  assign queue_bits_wb_pc__T_130_mask = 1'h0;
  assign queue_bits_wb_pc__T_130_en = reset;
  assign queue_bits_wb_pc__T_131_data = 32'h0;
  assign queue_bits_wb_pc__T_131_addr = 6'h3d;
  assign queue_bits_wb_pc__T_131_mask = 1'h0;
  assign queue_bits_wb_pc__T_131_en = reset;
  assign queue_bits_wb_pc__T_132_data = 32'h0;
  assign queue_bits_wb_pc__T_132_addr = 6'h3e;
  assign queue_bits_wb_pc__T_132_mask = 1'h0;
  assign queue_bits_wb_pc__T_132_en = reset;
  assign queue_bits_wb_pc__T_133_data = 32'h0;
  assign queue_bits_wb_pc__T_133_addr = 6'h3f;
  assign queue_bits_wb_pc__T_133_mask = 1'h0;
  assign queue_bits_wb_pc__T_133_en = reset;
  assign queue_bits_wb_pc_q_head_w_data = 32'h0;
  assign queue_bits_wb_pc_q_head_w_addr = head;
  assign queue_bits_wb_pc_q_head_w_mask = 1'h0;
  assign queue_bits_wb_pc_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_instr_op_q_head_r_addr = head;
  assign queue_bits_wb_instr_op_q_head_r_data = queue_bits_wb_instr_op[queue_bits_wb_instr_op_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_instr_op__T_3_data = io_enq_0_bits_data_wb_instr_op;
  assign queue_bits_wb_instr_op__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_instr_op__T_3_mask = 1'h1;
  assign queue_bits_wb_instr_op__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_instr_op__T_4_data = io_enq_1_bits_data_wb_instr_op;
  assign queue_bits_wb_instr_op__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_instr_op__T_4_mask = 1'h1;
  assign queue_bits_wb_instr_op__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_instr_op__T_5_data = 6'h0;
  assign queue_bits_wb_instr_op__T_5_addr = 6'h0;
  assign queue_bits_wb_instr_op__T_5_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_5_en = 1'h0;
  assign queue_bits_wb_instr_op__T_6_data = 6'h0;
  assign queue_bits_wb_instr_op__T_6_addr = 6'h1;
  assign queue_bits_wb_instr_op__T_6_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_6_en = 1'h0;
  assign queue_bits_wb_instr_op__T_7_data = 6'h0;
  assign queue_bits_wb_instr_op__T_7_addr = 6'h2;
  assign queue_bits_wb_instr_op__T_7_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_7_en = 1'h0;
  assign queue_bits_wb_instr_op__T_8_data = 6'h0;
  assign queue_bits_wb_instr_op__T_8_addr = 6'h3;
  assign queue_bits_wb_instr_op__T_8_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_8_en = 1'h0;
  assign queue_bits_wb_instr_op__T_9_data = 6'h0;
  assign queue_bits_wb_instr_op__T_9_addr = 6'h4;
  assign queue_bits_wb_instr_op__T_9_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_9_en = 1'h0;
  assign queue_bits_wb_instr_op__T_10_data = 6'h0;
  assign queue_bits_wb_instr_op__T_10_addr = 6'h5;
  assign queue_bits_wb_instr_op__T_10_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_10_en = 1'h0;
  assign queue_bits_wb_instr_op__T_11_data = 6'h0;
  assign queue_bits_wb_instr_op__T_11_addr = 6'h6;
  assign queue_bits_wb_instr_op__T_11_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_11_en = 1'h0;
  assign queue_bits_wb_instr_op__T_12_data = 6'h0;
  assign queue_bits_wb_instr_op__T_12_addr = 6'h7;
  assign queue_bits_wb_instr_op__T_12_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_12_en = 1'h0;
  assign queue_bits_wb_instr_op__T_13_data = 6'h0;
  assign queue_bits_wb_instr_op__T_13_addr = 6'h8;
  assign queue_bits_wb_instr_op__T_13_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_13_en = 1'h0;
  assign queue_bits_wb_instr_op__T_14_data = 6'h0;
  assign queue_bits_wb_instr_op__T_14_addr = 6'h9;
  assign queue_bits_wb_instr_op__T_14_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_14_en = 1'h0;
  assign queue_bits_wb_instr_op__T_15_data = 6'h0;
  assign queue_bits_wb_instr_op__T_15_addr = 6'ha;
  assign queue_bits_wb_instr_op__T_15_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_15_en = 1'h0;
  assign queue_bits_wb_instr_op__T_16_data = 6'h0;
  assign queue_bits_wb_instr_op__T_16_addr = 6'hb;
  assign queue_bits_wb_instr_op__T_16_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_16_en = 1'h0;
  assign queue_bits_wb_instr_op__T_17_data = 6'h0;
  assign queue_bits_wb_instr_op__T_17_addr = 6'hc;
  assign queue_bits_wb_instr_op__T_17_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_17_en = 1'h0;
  assign queue_bits_wb_instr_op__T_18_data = 6'h0;
  assign queue_bits_wb_instr_op__T_18_addr = 6'hd;
  assign queue_bits_wb_instr_op__T_18_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_18_en = 1'h0;
  assign queue_bits_wb_instr_op__T_19_data = 6'h0;
  assign queue_bits_wb_instr_op__T_19_addr = 6'he;
  assign queue_bits_wb_instr_op__T_19_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_19_en = 1'h0;
  assign queue_bits_wb_instr_op__T_20_data = 6'h0;
  assign queue_bits_wb_instr_op__T_20_addr = 6'hf;
  assign queue_bits_wb_instr_op__T_20_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_20_en = 1'h0;
  assign queue_bits_wb_instr_op__T_21_data = 6'h0;
  assign queue_bits_wb_instr_op__T_21_addr = 6'h10;
  assign queue_bits_wb_instr_op__T_21_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_21_en = 1'h0;
  assign queue_bits_wb_instr_op__T_22_data = 6'h0;
  assign queue_bits_wb_instr_op__T_22_addr = 6'h11;
  assign queue_bits_wb_instr_op__T_22_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_22_en = 1'h0;
  assign queue_bits_wb_instr_op__T_23_data = 6'h0;
  assign queue_bits_wb_instr_op__T_23_addr = 6'h12;
  assign queue_bits_wb_instr_op__T_23_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_23_en = 1'h0;
  assign queue_bits_wb_instr_op__T_24_data = 6'h0;
  assign queue_bits_wb_instr_op__T_24_addr = 6'h13;
  assign queue_bits_wb_instr_op__T_24_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_24_en = 1'h0;
  assign queue_bits_wb_instr_op__T_25_data = 6'h0;
  assign queue_bits_wb_instr_op__T_25_addr = 6'h14;
  assign queue_bits_wb_instr_op__T_25_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_25_en = 1'h0;
  assign queue_bits_wb_instr_op__T_26_data = 6'h0;
  assign queue_bits_wb_instr_op__T_26_addr = 6'h15;
  assign queue_bits_wb_instr_op__T_26_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_26_en = 1'h0;
  assign queue_bits_wb_instr_op__T_27_data = 6'h0;
  assign queue_bits_wb_instr_op__T_27_addr = 6'h16;
  assign queue_bits_wb_instr_op__T_27_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_27_en = 1'h0;
  assign queue_bits_wb_instr_op__T_28_data = 6'h0;
  assign queue_bits_wb_instr_op__T_28_addr = 6'h17;
  assign queue_bits_wb_instr_op__T_28_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_28_en = 1'h0;
  assign queue_bits_wb_instr_op__T_29_data = 6'h0;
  assign queue_bits_wb_instr_op__T_29_addr = 6'h18;
  assign queue_bits_wb_instr_op__T_29_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_29_en = 1'h0;
  assign queue_bits_wb_instr_op__T_30_data = 6'h0;
  assign queue_bits_wb_instr_op__T_30_addr = 6'h19;
  assign queue_bits_wb_instr_op__T_30_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_30_en = 1'h0;
  assign queue_bits_wb_instr_op__T_31_data = 6'h0;
  assign queue_bits_wb_instr_op__T_31_addr = 6'h1a;
  assign queue_bits_wb_instr_op__T_31_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_31_en = 1'h0;
  assign queue_bits_wb_instr_op__T_32_data = 6'h0;
  assign queue_bits_wb_instr_op__T_32_addr = 6'h1b;
  assign queue_bits_wb_instr_op__T_32_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_32_en = 1'h0;
  assign queue_bits_wb_instr_op__T_33_data = 6'h0;
  assign queue_bits_wb_instr_op__T_33_addr = 6'h1c;
  assign queue_bits_wb_instr_op__T_33_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_33_en = 1'h0;
  assign queue_bits_wb_instr_op__T_34_data = 6'h0;
  assign queue_bits_wb_instr_op__T_34_addr = 6'h1d;
  assign queue_bits_wb_instr_op__T_34_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_34_en = 1'h0;
  assign queue_bits_wb_instr_op__T_35_data = 6'h0;
  assign queue_bits_wb_instr_op__T_35_addr = 6'h1e;
  assign queue_bits_wb_instr_op__T_35_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_35_en = 1'h0;
  assign queue_bits_wb_instr_op__T_36_data = 6'h0;
  assign queue_bits_wb_instr_op__T_36_addr = 6'h1f;
  assign queue_bits_wb_instr_op__T_36_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_36_en = 1'h0;
  assign queue_bits_wb_instr_op__T_37_data = 6'h0;
  assign queue_bits_wb_instr_op__T_37_addr = 6'h20;
  assign queue_bits_wb_instr_op__T_37_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_37_en = 1'h0;
  assign queue_bits_wb_instr_op__T_38_data = 6'h0;
  assign queue_bits_wb_instr_op__T_38_addr = 6'h21;
  assign queue_bits_wb_instr_op__T_38_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_38_en = 1'h0;
  assign queue_bits_wb_instr_op__T_39_data = 6'h0;
  assign queue_bits_wb_instr_op__T_39_addr = 6'h22;
  assign queue_bits_wb_instr_op__T_39_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_39_en = 1'h0;
  assign queue_bits_wb_instr_op__T_40_data = 6'h0;
  assign queue_bits_wb_instr_op__T_40_addr = 6'h23;
  assign queue_bits_wb_instr_op__T_40_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_40_en = 1'h0;
  assign queue_bits_wb_instr_op__T_41_data = 6'h0;
  assign queue_bits_wb_instr_op__T_41_addr = 6'h24;
  assign queue_bits_wb_instr_op__T_41_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_41_en = 1'h0;
  assign queue_bits_wb_instr_op__T_42_data = 6'h0;
  assign queue_bits_wb_instr_op__T_42_addr = 6'h25;
  assign queue_bits_wb_instr_op__T_42_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_42_en = 1'h0;
  assign queue_bits_wb_instr_op__T_43_data = 6'h0;
  assign queue_bits_wb_instr_op__T_43_addr = 6'h26;
  assign queue_bits_wb_instr_op__T_43_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_43_en = 1'h0;
  assign queue_bits_wb_instr_op__T_44_data = 6'h0;
  assign queue_bits_wb_instr_op__T_44_addr = 6'h27;
  assign queue_bits_wb_instr_op__T_44_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_44_en = 1'h0;
  assign queue_bits_wb_instr_op__T_45_data = 6'h0;
  assign queue_bits_wb_instr_op__T_45_addr = 6'h28;
  assign queue_bits_wb_instr_op__T_45_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_45_en = 1'h0;
  assign queue_bits_wb_instr_op__T_46_data = 6'h0;
  assign queue_bits_wb_instr_op__T_46_addr = 6'h29;
  assign queue_bits_wb_instr_op__T_46_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_46_en = 1'h0;
  assign queue_bits_wb_instr_op__T_47_data = 6'h0;
  assign queue_bits_wb_instr_op__T_47_addr = 6'h2a;
  assign queue_bits_wb_instr_op__T_47_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_47_en = 1'h0;
  assign queue_bits_wb_instr_op__T_48_data = 6'h0;
  assign queue_bits_wb_instr_op__T_48_addr = 6'h2b;
  assign queue_bits_wb_instr_op__T_48_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_48_en = 1'h0;
  assign queue_bits_wb_instr_op__T_49_data = 6'h0;
  assign queue_bits_wb_instr_op__T_49_addr = 6'h2c;
  assign queue_bits_wb_instr_op__T_49_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_49_en = 1'h0;
  assign queue_bits_wb_instr_op__T_50_data = 6'h0;
  assign queue_bits_wb_instr_op__T_50_addr = 6'h2d;
  assign queue_bits_wb_instr_op__T_50_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_50_en = 1'h0;
  assign queue_bits_wb_instr_op__T_51_data = 6'h0;
  assign queue_bits_wb_instr_op__T_51_addr = 6'h2e;
  assign queue_bits_wb_instr_op__T_51_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_51_en = 1'h0;
  assign queue_bits_wb_instr_op__T_52_data = 6'h0;
  assign queue_bits_wb_instr_op__T_52_addr = 6'h2f;
  assign queue_bits_wb_instr_op__T_52_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_52_en = 1'h0;
  assign queue_bits_wb_instr_op__T_53_data = 6'h0;
  assign queue_bits_wb_instr_op__T_53_addr = 6'h30;
  assign queue_bits_wb_instr_op__T_53_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_53_en = 1'h0;
  assign queue_bits_wb_instr_op__T_54_data = 6'h0;
  assign queue_bits_wb_instr_op__T_54_addr = 6'h31;
  assign queue_bits_wb_instr_op__T_54_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_54_en = 1'h0;
  assign queue_bits_wb_instr_op__T_55_data = 6'h0;
  assign queue_bits_wb_instr_op__T_55_addr = 6'h32;
  assign queue_bits_wb_instr_op__T_55_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_55_en = 1'h0;
  assign queue_bits_wb_instr_op__T_56_data = 6'h0;
  assign queue_bits_wb_instr_op__T_56_addr = 6'h33;
  assign queue_bits_wb_instr_op__T_56_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_56_en = 1'h0;
  assign queue_bits_wb_instr_op__T_57_data = 6'h0;
  assign queue_bits_wb_instr_op__T_57_addr = 6'h34;
  assign queue_bits_wb_instr_op__T_57_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_57_en = 1'h0;
  assign queue_bits_wb_instr_op__T_58_data = 6'h0;
  assign queue_bits_wb_instr_op__T_58_addr = 6'h35;
  assign queue_bits_wb_instr_op__T_58_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_58_en = 1'h0;
  assign queue_bits_wb_instr_op__T_59_data = 6'h0;
  assign queue_bits_wb_instr_op__T_59_addr = 6'h36;
  assign queue_bits_wb_instr_op__T_59_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_59_en = 1'h0;
  assign queue_bits_wb_instr_op__T_60_data = 6'h0;
  assign queue_bits_wb_instr_op__T_60_addr = 6'h37;
  assign queue_bits_wb_instr_op__T_60_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_60_en = 1'h0;
  assign queue_bits_wb_instr_op__T_61_data = 6'h0;
  assign queue_bits_wb_instr_op__T_61_addr = 6'h38;
  assign queue_bits_wb_instr_op__T_61_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_61_en = 1'h0;
  assign queue_bits_wb_instr_op__T_62_data = 6'h0;
  assign queue_bits_wb_instr_op__T_62_addr = 6'h39;
  assign queue_bits_wb_instr_op__T_62_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_62_en = 1'h0;
  assign queue_bits_wb_instr_op__T_63_data = 6'h0;
  assign queue_bits_wb_instr_op__T_63_addr = 6'h3a;
  assign queue_bits_wb_instr_op__T_63_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_63_en = 1'h0;
  assign queue_bits_wb_instr_op__T_64_data = 6'h0;
  assign queue_bits_wb_instr_op__T_64_addr = 6'h3b;
  assign queue_bits_wb_instr_op__T_64_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_64_en = 1'h0;
  assign queue_bits_wb_instr_op__T_65_data = 6'h0;
  assign queue_bits_wb_instr_op__T_65_addr = 6'h3c;
  assign queue_bits_wb_instr_op__T_65_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_65_en = 1'h0;
  assign queue_bits_wb_instr_op__T_66_data = 6'h0;
  assign queue_bits_wb_instr_op__T_66_addr = 6'h3d;
  assign queue_bits_wb_instr_op__T_66_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_66_en = 1'h0;
  assign queue_bits_wb_instr_op__T_67_data = 6'h0;
  assign queue_bits_wb_instr_op__T_67_addr = 6'h3e;
  assign queue_bits_wb_instr_op__T_67_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_67_en = 1'h0;
  assign queue_bits_wb_instr_op__T_68_data = 6'h0;
  assign queue_bits_wb_instr_op__T_68_addr = 6'h3f;
  assign queue_bits_wb_instr_op__T_68_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_68_en = 1'h0;
  assign queue_bits_wb_instr_op__T_70_data = 6'h0;
  assign queue_bits_wb_instr_op__T_70_addr = 6'h0;
  assign queue_bits_wb_instr_op__T_70_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_70_en = reset;
  assign queue_bits_wb_instr_op__T_71_data = 6'h0;
  assign queue_bits_wb_instr_op__T_71_addr = 6'h1;
  assign queue_bits_wb_instr_op__T_71_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_71_en = reset;
  assign queue_bits_wb_instr_op__T_72_data = 6'h0;
  assign queue_bits_wb_instr_op__T_72_addr = 6'h2;
  assign queue_bits_wb_instr_op__T_72_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_72_en = reset;
  assign queue_bits_wb_instr_op__T_73_data = 6'h0;
  assign queue_bits_wb_instr_op__T_73_addr = 6'h3;
  assign queue_bits_wb_instr_op__T_73_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_73_en = reset;
  assign queue_bits_wb_instr_op__T_74_data = 6'h0;
  assign queue_bits_wb_instr_op__T_74_addr = 6'h4;
  assign queue_bits_wb_instr_op__T_74_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_74_en = reset;
  assign queue_bits_wb_instr_op__T_75_data = 6'h0;
  assign queue_bits_wb_instr_op__T_75_addr = 6'h5;
  assign queue_bits_wb_instr_op__T_75_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_75_en = reset;
  assign queue_bits_wb_instr_op__T_76_data = 6'h0;
  assign queue_bits_wb_instr_op__T_76_addr = 6'h6;
  assign queue_bits_wb_instr_op__T_76_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_76_en = reset;
  assign queue_bits_wb_instr_op__T_77_data = 6'h0;
  assign queue_bits_wb_instr_op__T_77_addr = 6'h7;
  assign queue_bits_wb_instr_op__T_77_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_77_en = reset;
  assign queue_bits_wb_instr_op__T_78_data = 6'h0;
  assign queue_bits_wb_instr_op__T_78_addr = 6'h8;
  assign queue_bits_wb_instr_op__T_78_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_78_en = reset;
  assign queue_bits_wb_instr_op__T_79_data = 6'h0;
  assign queue_bits_wb_instr_op__T_79_addr = 6'h9;
  assign queue_bits_wb_instr_op__T_79_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_79_en = reset;
  assign queue_bits_wb_instr_op__T_80_data = 6'h0;
  assign queue_bits_wb_instr_op__T_80_addr = 6'ha;
  assign queue_bits_wb_instr_op__T_80_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_80_en = reset;
  assign queue_bits_wb_instr_op__T_81_data = 6'h0;
  assign queue_bits_wb_instr_op__T_81_addr = 6'hb;
  assign queue_bits_wb_instr_op__T_81_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_81_en = reset;
  assign queue_bits_wb_instr_op__T_82_data = 6'h0;
  assign queue_bits_wb_instr_op__T_82_addr = 6'hc;
  assign queue_bits_wb_instr_op__T_82_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_82_en = reset;
  assign queue_bits_wb_instr_op__T_83_data = 6'h0;
  assign queue_bits_wb_instr_op__T_83_addr = 6'hd;
  assign queue_bits_wb_instr_op__T_83_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_83_en = reset;
  assign queue_bits_wb_instr_op__T_84_data = 6'h0;
  assign queue_bits_wb_instr_op__T_84_addr = 6'he;
  assign queue_bits_wb_instr_op__T_84_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_84_en = reset;
  assign queue_bits_wb_instr_op__T_85_data = 6'h0;
  assign queue_bits_wb_instr_op__T_85_addr = 6'hf;
  assign queue_bits_wb_instr_op__T_85_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_85_en = reset;
  assign queue_bits_wb_instr_op__T_86_data = 6'h0;
  assign queue_bits_wb_instr_op__T_86_addr = 6'h10;
  assign queue_bits_wb_instr_op__T_86_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_86_en = reset;
  assign queue_bits_wb_instr_op__T_87_data = 6'h0;
  assign queue_bits_wb_instr_op__T_87_addr = 6'h11;
  assign queue_bits_wb_instr_op__T_87_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_87_en = reset;
  assign queue_bits_wb_instr_op__T_88_data = 6'h0;
  assign queue_bits_wb_instr_op__T_88_addr = 6'h12;
  assign queue_bits_wb_instr_op__T_88_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_88_en = reset;
  assign queue_bits_wb_instr_op__T_89_data = 6'h0;
  assign queue_bits_wb_instr_op__T_89_addr = 6'h13;
  assign queue_bits_wb_instr_op__T_89_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_89_en = reset;
  assign queue_bits_wb_instr_op__T_90_data = 6'h0;
  assign queue_bits_wb_instr_op__T_90_addr = 6'h14;
  assign queue_bits_wb_instr_op__T_90_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_90_en = reset;
  assign queue_bits_wb_instr_op__T_91_data = 6'h0;
  assign queue_bits_wb_instr_op__T_91_addr = 6'h15;
  assign queue_bits_wb_instr_op__T_91_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_91_en = reset;
  assign queue_bits_wb_instr_op__T_92_data = 6'h0;
  assign queue_bits_wb_instr_op__T_92_addr = 6'h16;
  assign queue_bits_wb_instr_op__T_92_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_92_en = reset;
  assign queue_bits_wb_instr_op__T_93_data = 6'h0;
  assign queue_bits_wb_instr_op__T_93_addr = 6'h17;
  assign queue_bits_wb_instr_op__T_93_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_93_en = reset;
  assign queue_bits_wb_instr_op__T_94_data = 6'h0;
  assign queue_bits_wb_instr_op__T_94_addr = 6'h18;
  assign queue_bits_wb_instr_op__T_94_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_94_en = reset;
  assign queue_bits_wb_instr_op__T_95_data = 6'h0;
  assign queue_bits_wb_instr_op__T_95_addr = 6'h19;
  assign queue_bits_wb_instr_op__T_95_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_95_en = reset;
  assign queue_bits_wb_instr_op__T_96_data = 6'h0;
  assign queue_bits_wb_instr_op__T_96_addr = 6'h1a;
  assign queue_bits_wb_instr_op__T_96_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_96_en = reset;
  assign queue_bits_wb_instr_op__T_97_data = 6'h0;
  assign queue_bits_wb_instr_op__T_97_addr = 6'h1b;
  assign queue_bits_wb_instr_op__T_97_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_97_en = reset;
  assign queue_bits_wb_instr_op__T_98_data = 6'h0;
  assign queue_bits_wb_instr_op__T_98_addr = 6'h1c;
  assign queue_bits_wb_instr_op__T_98_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_98_en = reset;
  assign queue_bits_wb_instr_op__T_99_data = 6'h0;
  assign queue_bits_wb_instr_op__T_99_addr = 6'h1d;
  assign queue_bits_wb_instr_op__T_99_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_99_en = reset;
  assign queue_bits_wb_instr_op__T_100_data = 6'h0;
  assign queue_bits_wb_instr_op__T_100_addr = 6'h1e;
  assign queue_bits_wb_instr_op__T_100_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_100_en = reset;
  assign queue_bits_wb_instr_op__T_101_data = 6'h0;
  assign queue_bits_wb_instr_op__T_101_addr = 6'h1f;
  assign queue_bits_wb_instr_op__T_101_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_101_en = reset;
  assign queue_bits_wb_instr_op__T_102_data = 6'h0;
  assign queue_bits_wb_instr_op__T_102_addr = 6'h20;
  assign queue_bits_wb_instr_op__T_102_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_102_en = reset;
  assign queue_bits_wb_instr_op__T_103_data = 6'h0;
  assign queue_bits_wb_instr_op__T_103_addr = 6'h21;
  assign queue_bits_wb_instr_op__T_103_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_103_en = reset;
  assign queue_bits_wb_instr_op__T_104_data = 6'h0;
  assign queue_bits_wb_instr_op__T_104_addr = 6'h22;
  assign queue_bits_wb_instr_op__T_104_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_104_en = reset;
  assign queue_bits_wb_instr_op__T_105_data = 6'h0;
  assign queue_bits_wb_instr_op__T_105_addr = 6'h23;
  assign queue_bits_wb_instr_op__T_105_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_105_en = reset;
  assign queue_bits_wb_instr_op__T_106_data = 6'h0;
  assign queue_bits_wb_instr_op__T_106_addr = 6'h24;
  assign queue_bits_wb_instr_op__T_106_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_106_en = reset;
  assign queue_bits_wb_instr_op__T_107_data = 6'h0;
  assign queue_bits_wb_instr_op__T_107_addr = 6'h25;
  assign queue_bits_wb_instr_op__T_107_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_107_en = reset;
  assign queue_bits_wb_instr_op__T_108_data = 6'h0;
  assign queue_bits_wb_instr_op__T_108_addr = 6'h26;
  assign queue_bits_wb_instr_op__T_108_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_108_en = reset;
  assign queue_bits_wb_instr_op__T_109_data = 6'h0;
  assign queue_bits_wb_instr_op__T_109_addr = 6'h27;
  assign queue_bits_wb_instr_op__T_109_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_109_en = reset;
  assign queue_bits_wb_instr_op__T_110_data = 6'h0;
  assign queue_bits_wb_instr_op__T_110_addr = 6'h28;
  assign queue_bits_wb_instr_op__T_110_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_110_en = reset;
  assign queue_bits_wb_instr_op__T_111_data = 6'h0;
  assign queue_bits_wb_instr_op__T_111_addr = 6'h29;
  assign queue_bits_wb_instr_op__T_111_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_111_en = reset;
  assign queue_bits_wb_instr_op__T_112_data = 6'h0;
  assign queue_bits_wb_instr_op__T_112_addr = 6'h2a;
  assign queue_bits_wb_instr_op__T_112_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_112_en = reset;
  assign queue_bits_wb_instr_op__T_113_data = 6'h0;
  assign queue_bits_wb_instr_op__T_113_addr = 6'h2b;
  assign queue_bits_wb_instr_op__T_113_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_113_en = reset;
  assign queue_bits_wb_instr_op__T_114_data = 6'h0;
  assign queue_bits_wb_instr_op__T_114_addr = 6'h2c;
  assign queue_bits_wb_instr_op__T_114_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_114_en = reset;
  assign queue_bits_wb_instr_op__T_115_data = 6'h0;
  assign queue_bits_wb_instr_op__T_115_addr = 6'h2d;
  assign queue_bits_wb_instr_op__T_115_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_115_en = reset;
  assign queue_bits_wb_instr_op__T_116_data = 6'h0;
  assign queue_bits_wb_instr_op__T_116_addr = 6'h2e;
  assign queue_bits_wb_instr_op__T_116_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_116_en = reset;
  assign queue_bits_wb_instr_op__T_117_data = 6'h0;
  assign queue_bits_wb_instr_op__T_117_addr = 6'h2f;
  assign queue_bits_wb_instr_op__T_117_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_117_en = reset;
  assign queue_bits_wb_instr_op__T_118_data = 6'h0;
  assign queue_bits_wb_instr_op__T_118_addr = 6'h30;
  assign queue_bits_wb_instr_op__T_118_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_118_en = reset;
  assign queue_bits_wb_instr_op__T_119_data = 6'h0;
  assign queue_bits_wb_instr_op__T_119_addr = 6'h31;
  assign queue_bits_wb_instr_op__T_119_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_119_en = reset;
  assign queue_bits_wb_instr_op__T_120_data = 6'h0;
  assign queue_bits_wb_instr_op__T_120_addr = 6'h32;
  assign queue_bits_wb_instr_op__T_120_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_120_en = reset;
  assign queue_bits_wb_instr_op__T_121_data = 6'h0;
  assign queue_bits_wb_instr_op__T_121_addr = 6'h33;
  assign queue_bits_wb_instr_op__T_121_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_121_en = reset;
  assign queue_bits_wb_instr_op__T_122_data = 6'h0;
  assign queue_bits_wb_instr_op__T_122_addr = 6'h34;
  assign queue_bits_wb_instr_op__T_122_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_122_en = reset;
  assign queue_bits_wb_instr_op__T_123_data = 6'h0;
  assign queue_bits_wb_instr_op__T_123_addr = 6'h35;
  assign queue_bits_wb_instr_op__T_123_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_123_en = reset;
  assign queue_bits_wb_instr_op__T_124_data = 6'h0;
  assign queue_bits_wb_instr_op__T_124_addr = 6'h36;
  assign queue_bits_wb_instr_op__T_124_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_124_en = reset;
  assign queue_bits_wb_instr_op__T_125_data = 6'h0;
  assign queue_bits_wb_instr_op__T_125_addr = 6'h37;
  assign queue_bits_wb_instr_op__T_125_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_125_en = reset;
  assign queue_bits_wb_instr_op__T_126_data = 6'h0;
  assign queue_bits_wb_instr_op__T_126_addr = 6'h38;
  assign queue_bits_wb_instr_op__T_126_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_126_en = reset;
  assign queue_bits_wb_instr_op__T_127_data = 6'h0;
  assign queue_bits_wb_instr_op__T_127_addr = 6'h39;
  assign queue_bits_wb_instr_op__T_127_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_127_en = reset;
  assign queue_bits_wb_instr_op__T_128_data = 6'h0;
  assign queue_bits_wb_instr_op__T_128_addr = 6'h3a;
  assign queue_bits_wb_instr_op__T_128_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_128_en = reset;
  assign queue_bits_wb_instr_op__T_129_data = 6'h0;
  assign queue_bits_wb_instr_op__T_129_addr = 6'h3b;
  assign queue_bits_wb_instr_op__T_129_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_129_en = reset;
  assign queue_bits_wb_instr_op__T_130_data = 6'h0;
  assign queue_bits_wb_instr_op__T_130_addr = 6'h3c;
  assign queue_bits_wb_instr_op__T_130_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_130_en = reset;
  assign queue_bits_wb_instr_op__T_131_data = 6'h0;
  assign queue_bits_wb_instr_op__T_131_addr = 6'h3d;
  assign queue_bits_wb_instr_op__T_131_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_131_en = reset;
  assign queue_bits_wb_instr_op__T_132_data = 6'h0;
  assign queue_bits_wb_instr_op__T_132_addr = 6'h3e;
  assign queue_bits_wb_instr_op__T_132_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_132_en = reset;
  assign queue_bits_wb_instr_op__T_133_data = 6'h0;
  assign queue_bits_wb_instr_op__T_133_addr = 6'h3f;
  assign queue_bits_wb_instr_op__T_133_mask = 1'h0;
  assign queue_bits_wb_instr_op__T_133_en = reset;
  assign queue_bits_wb_instr_op_q_head_w_data = 6'h0;
  assign queue_bits_wb_instr_op_q_head_w_addr = head;
  assign queue_bits_wb_instr_op_q_head_w_mask = 1'h0;
  assign queue_bits_wb_instr_op_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_instr_rs_idx_q_head_r_addr = head;
  assign queue_bits_wb_instr_rs_idx_q_head_r_data = queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_instr_rs_idx__T_3_data = io_enq_0_bits_data_wb_instr_rs_idx;
  assign queue_bits_wb_instr_rs_idx__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_instr_rs_idx__T_3_mask = 1'h1;
  assign queue_bits_wb_instr_rs_idx__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_instr_rs_idx__T_4_data = io_enq_1_bits_data_wb_instr_rs_idx;
  assign queue_bits_wb_instr_rs_idx__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_instr_rs_idx__T_4_mask = 1'h1;
  assign queue_bits_wb_instr_rs_idx__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_instr_rs_idx__T_5_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_5_addr = 6'h0;
  assign queue_bits_wb_instr_rs_idx__T_5_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_5_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_6_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_6_addr = 6'h1;
  assign queue_bits_wb_instr_rs_idx__T_6_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_6_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_7_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_7_addr = 6'h2;
  assign queue_bits_wb_instr_rs_idx__T_7_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_7_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_8_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_8_addr = 6'h3;
  assign queue_bits_wb_instr_rs_idx__T_8_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_8_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_9_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_9_addr = 6'h4;
  assign queue_bits_wb_instr_rs_idx__T_9_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_9_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_10_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_10_addr = 6'h5;
  assign queue_bits_wb_instr_rs_idx__T_10_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_10_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_11_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_11_addr = 6'h6;
  assign queue_bits_wb_instr_rs_idx__T_11_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_11_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_12_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_12_addr = 6'h7;
  assign queue_bits_wb_instr_rs_idx__T_12_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_12_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_13_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_13_addr = 6'h8;
  assign queue_bits_wb_instr_rs_idx__T_13_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_13_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_14_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_14_addr = 6'h9;
  assign queue_bits_wb_instr_rs_idx__T_14_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_14_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_15_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_15_addr = 6'ha;
  assign queue_bits_wb_instr_rs_idx__T_15_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_15_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_16_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_16_addr = 6'hb;
  assign queue_bits_wb_instr_rs_idx__T_16_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_16_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_17_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_17_addr = 6'hc;
  assign queue_bits_wb_instr_rs_idx__T_17_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_17_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_18_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_18_addr = 6'hd;
  assign queue_bits_wb_instr_rs_idx__T_18_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_18_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_19_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_19_addr = 6'he;
  assign queue_bits_wb_instr_rs_idx__T_19_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_19_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_20_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_20_addr = 6'hf;
  assign queue_bits_wb_instr_rs_idx__T_20_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_20_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_21_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_21_addr = 6'h10;
  assign queue_bits_wb_instr_rs_idx__T_21_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_21_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_22_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_22_addr = 6'h11;
  assign queue_bits_wb_instr_rs_idx__T_22_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_22_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_23_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_23_addr = 6'h12;
  assign queue_bits_wb_instr_rs_idx__T_23_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_23_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_24_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_24_addr = 6'h13;
  assign queue_bits_wb_instr_rs_idx__T_24_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_24_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_25_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_25_addr = 6'h14;
  assign queue_bits_wb_instr_rs_idx__T_25_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_25_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_26_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_26_addr = 6'h15;
  assign queue_bits_wb_instr_rs_idx__T_26_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_26_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_27_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_27_addr = 6'h16;
  assign queue_bits_wb_instr_rs_idx__T_27_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_27_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_28_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_28_addr = 6'h17;
  assign queue_bits_wb_instr_rs_idx__T_28_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_28_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_29_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_29_addr = 6'h18;
  assign queue_bits_wb_instr_rs_idx__T_29_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_29_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_30_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_30_addr = 6'h19;
  assign queue_bits_wb_instr_rs_idx__T_30_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_30_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_31_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_31_addr = 6'h1a;
  assign queue_bits_wb_instr_rs_idx__T_31_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_31_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_32_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_32_addr = 6'h1b;
  assign queue_bits_wb_instr_rs_idx__T_32_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_32_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_33_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_33_addr = 6'h1c;
  assign queue_bits_wb_instr_rs_idx__T_33_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_33_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_34_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_34_addr = 6'h1d;
  assign queue_bits_wb_instr_rs_idx__T_34_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_34_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_35_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_35_addr = 6'h1e;
  assign queue_bits_wb_instr_rs_idx__T_35_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_35_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_36_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_36_addr = 6'h1f;
  assign queue_bits_wb_instr_rs_idx__T_36_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_36_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_37_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_37_addr = 6'h20;
  assign queue_bits_wb_instr_rs_idx__T_37_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_37_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_38_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_38_addr = 6'h21;
  assign queue_bits_wb_instr_rs_idx__T_38_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_38_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_39_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_39_addr = 6'h22;
  assign queue_bits_wb_instr_rs_idx__T_39_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_39_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_40_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_40_addr = 6'h23;
  assign queue_bits_wb_instr_rs_idx__T_40_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_40_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_41_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_41_addr = 6'h24;
  assign queue_bits_wb_instr_rs_idx__T_41_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_41_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_42_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_42_addr = 6'h25;
  assign queue_bits_wb_instr_rs_idx__T_42_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_42_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_43_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_43_addr = 6'h26;
  assign queue_bits_wb_instr_rs_idx__T_43_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_43_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_44_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_44_addr = 6'h27;
  assign queue_bits_wb_instr_rs_idx__T_44_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_44_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_45_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_45_addr = 6'h28;
  assign queue_bits_wb_instr_rs_idx__T_45_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_45_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_46_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_46_addr = 6'h29;
  assign queue_bits_wb_instr_rs_idx__T_46_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_46_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_47_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_47_addr = 6'h2a;
  assign queue_bits_wb_instr_rs_idx__T_47_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_47_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_48_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_48_addr = 6'h2b;
  assign queue_bits_wb_instr_rs_idx__T_48_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_48_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_49_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_49_addr = 6'h2c;
  assign queue_bits_wb_instr_rs_idx__T_49_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_49_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_50_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_50_addr = 6'h2d;
  assign queue_bits_wb_instr_rs_idx__T_50_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_50_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_51_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_51_addr = 6'h2e;
  assign queue_bits_wb_instr_rs_idx__T_51_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_51_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_52_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_52_addr = 6'h2f;
  assign queue_bits_wb_instr_rs_idx__T_52_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_52_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_53_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_53_addr = 6'h30;
  assign queue_bits_wb_instr_rs_idx__T_53_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_53_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_54_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_54_addr = 6'h31;
  assign queue_bits_wb_instr_rs_idx__T_54_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_54_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_55_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_55_addr = 6'h32;
  assign queue_bits_wb_instr_rs_idx__T_55_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_55_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_56_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_56_addr = 6'h33;
  assign queue_bits_wb_instr_rs_idx__T_56_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_56_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_57_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_57_addr = 6'h34;
  assign queue_bits_wb_instr_rs_idx__T_57_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_57_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_58_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_58_addr = 6'h35;
  assign queue_bits_wb_instr_rs_idx__T_58_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_58_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_59_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_59_addr = 6'h36;
  assign queue_bits_wb_instr_rs_idx__T_59_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_59_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_60_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_60_addr = 6'h37;
  assign queue_bits_wb_instr_rs_idx__T_60_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_60_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_61_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_61_addr = 6'h38;
  assign queue_bits_wb_instr_rs_idx__T_61_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_61_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_62_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_62_addr = 6'h39;
  assign queue_bits_wb_instr_rs_idx__T_62_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_62_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_63_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_63_addr = 6'h3a;
  assign queue_bits_wb_instr_rs_idx__T_63_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_63_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_64_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_64_addr = 6'h3b;
  assign queue_bits_wb_instr_rs_idx__T_64_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_64_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_65_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_65_addr = 6'h3c;
  assign queue_bits_wb_instr_rs_idx__T_65_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_65_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_66_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_66_addr = 6'h3d;
  assign queue_bits_wb_instr_rs_idx__T_66_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_66_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_67_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_67_addr = 6'h3e;
  assign queue_bits_wb_instr_rs_idx__T_67_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_67_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_68_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_68_addr = 6'h3f;
  assign queue_bits_wb_instr_rs_idx__T_68_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_68_en = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_70_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_70_addr = 6'h0;
  assign queue_bits_wb_instr_rs_idx__T_70_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_70_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_71_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_71_addr = 6'h1;
  assign queue_bits_wb_instr_rs_idx__T_71_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_71_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_72_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_72_addr = 6'h2;
  assign queue_bits_wb_instr_rs_idx__T_72_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_72_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_73_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_73_addr = 6'h3;
  assign queue_bits_wb_instr_rs_idx__T_73_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_73_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_74_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_74_addr = 6'h4;
  assign queue_bits_wb_instr_rs_idx__T_74_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_74_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_75_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_75_addr = 6'h5;
  assign queue_bits_wb_instr_rs_idx__T_75_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_75_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_76_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_76_addr = 6'h6;
  assign queue_bits_wb_instr_rs_idx__T_76_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_76_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_77_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_77_addr = 6'h7;
  assign queue_bits_wb_instr_rs_idx__T_77_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_77_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_78_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_78_addr = 6'h8;
  assign queue_bits_wb_instr_rs_idx__T_78_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_78_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_79_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_79_addr = 6'h9;
  assign queue_bits_wb_instr_rs_idx__T_79_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_79_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_80_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_80_addr = 6'ha;
  assign queue_bits_wb_instr_rs_idx__T_80_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_80_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_81_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_81_addr = 6'hb;
  assign queue_bits_wb_instr_rs_idx__T_81_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_81_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_82_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_82_addr = 6'hc;
  assign queue_bits_wb_instr_rs_idx__T_82_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_82_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_83_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_83_addr = 6'hd;
  assign queue_bits_wb_instr_rs_idx__T_83_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_83_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_84_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_84_addr = 6'he;
  assign queue_bits_wb_instr_rs_idx__T_84_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_84_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_85_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_85_addr = 6'hf;
  assign queue_bits_wb_instr_rs_idx__T_85_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_85_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_86_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_86_addr = 6'h10;
  assign queue_bits_wb_instr_rs_idx__T_86_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_86_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_87_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_87_addr = 6'h11;
  assign queue_bits_wb_instr_rs_idx__T_87_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_87_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_88_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_88_addr = 6'h12;
  assign queue_bits_wb_instr_rs_idx__T_88_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_88_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_89_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_89_addr = 6'h13;
  assign queue_bits_wb_instr_rs_idx__T_89_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_89_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_90_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_90_addr = 6'h14;
  assign queue_bits_wb_instr_rs_idx__T_90_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_90_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_91_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_91_addr = 6'h15;
  assign queue_bits_wb_instr_rs_idx__T_91_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_91_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_92_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_92_addr = 6'h16;
  assign queue_bits_wb_instr_rs_idx__T_92_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_92_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_93_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_93_addr = 6'h17;
  assign queue_bits_wb_instr_rs_idx__T_93_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_93_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_94_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_94_addr = 6'h18;
  assign queue_bits_wb_instr_rs_idx__T_94_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_94_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_95_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_95_addr = 6'h19;
  assign queue_bits_wb_instr_rs_idx__T_95_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_95_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_96_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_96_addr = 6'h1a;
  assign queue_bits_wb_instr_rs_idx__T_96_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_96_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_97_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_97_addr = 6'h1b;
  assign queue_bits_wb_instr_rs_idx__T_97_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_97_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_98_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_98_addr = 6'h1c;
  assign queue_bits_wb_instr_rs_idx__T_98_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_98_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_99_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_99_addr = 6'h1d;
  assign queue_bits_wb_instr_rs_idx__T_99_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_99_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_100_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_100_addr = 6'h1e;
  assign queue_bits_wb_instr_rs_idx__T_100_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_100_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_101_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_101_addr = 6'h1f;
  assign queue_bits_wb_instr_rs_idx__T_101_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_101_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_102_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_102_addr = 6'h20;
  assign queue_bits_wb_instr_rs_idx__T_102_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_102_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_103_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_103_addr = 6'h21;
  assign queue_bits_wb_instr_rs_idx__T_103_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_103_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_104_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_104_addr = 6'h22;
  assign queue_bits_wb_instr_rs_idx__T_104_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_104_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_105_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_105_addr = 6'h23;
  assign queue_bits_wb_instr_rs_idx__T_105_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_105_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_106_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_106_addr = 6'h24;
  assign queue_bits_wb_instr_rs_idx__T_106_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_106_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_107_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_107_addr = 6'h25;
  assign queue_bits_wb_instr_rs_idx__T_107_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_107_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_108_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_108_addr = 6'h26;
  assign queue_bits_wb_instr_rs_idx__T_108_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_108_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_109_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_109_addr = 6'h27;
  assign queue_bits_wb_instr_rs_idx__T_109_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_109_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_110_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_110_addr = 6'h28;
  assign queue_bits_wb_instr_rs_idx__T_110_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_110_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_111_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_111_addr = 6'h29;
  assign queue_bits_wb_instr_rs_idx__T_111_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_111_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_112_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_112_addr = 6'h2a;
  assign queue_bits_wb_instr_rs_idx__T_112_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_112_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_113_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_113_addr = 6'h2b;
  assign queue_bits_wb_instr_rs_idx__T_113_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_113_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_114_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_114_addr = 6'h2c;
  assign queue_bits_wb_instr_rs_idx__T_114_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_114_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_115_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_115_addr = 6'h2d;
  assign queue_bits_wb_instr_rs_idx__T_115_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_115_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_116_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_116_addr = 6'h2e;
  assign queue_bits_wb_instr_rs_idx__T_116_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_116_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_117_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_117_addr = 6'h2f;
  assign queue_bits_wb_instr_rs_idx__T_117_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_117_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_118_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_118_addr = 6'h30;
  assign queue_bits_wb_instr_rs_idx__T_118_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_118_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_119_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_119_addr = 6'h31;
  assign queue_bits_wb_instr_rs_idx__T_119_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_119_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_120_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_120_addr = 6'h32;
  assign queue_bits_wb_instr_rs_idx__T_120_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_120_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_121_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_121_addr = 6'h33;
  assign queue_bits_wb_instr_rs_idx__T_121_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_121_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_122_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_122_addr = 6'h34;
  assign queue_bits_wb_instr_rs_idx__T_122_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_122_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_123_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_123_addr = 6'h35;
  assign queue_bits_wb_instr_rs_idx__T_123_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_123_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_124_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_124_addr = 6'h36;
  assign queue_bits_wb_instr_rs_idx__T_124_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_124_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_125_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_125_addr = 6'h37;
  assign queue_bits_wb_instr_rs_idx__T_125_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_125_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_126_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_126_addr = 6'h38;
  assign queue_bits_wb_instr_rs_idx__T_126_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_126_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_127_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_127_addr = 6'h39;
  assign queue_bits_wb_instr_rs_idx__T_127_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_127_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_128_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_128_addr = 6'h3a;
  assign queue_bits_wb_instr_rs_idx__T_128_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_128_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_129_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_129_addr = 6'h3b;
  assign queue_bits_wb_instr_rs_idx__T_129_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_129_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_130_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_130_addr = 6'h3c;
  assign queue_bits_wb_instr_rs_idx__T_130_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_130_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_131_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_131_addr = 6'h3d;
  assign queue_bits_wb_instr_rs_idx__T_131_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_131_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_132_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_132_addr = 6'h3e;
  assign queue_bits_wb_instr_rs_idx__T_132_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_132_en = reset;
  assign queue_bits_wb_instr_rs_idx__T_133_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx__T_133_addr = 6'h3f;
  assign queue_bits_wb_instr_rs_idx__T_133_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx__T_133_en = reset;
  assign queue_bits_wb_instr_rs_idx_q_head_w_data = 5'h0;
  assign queue_bits_wb_instr_rs_idx_q_head_w_addr = head;
  assign queue_bits_wb_instr_rs_idx_q_head_w_mask = 1'h0;
  assign queue_bits_wb_instr_rs_idx_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_instr_rt_idx_q_head_r_addr = head;
  assign queue_bits_wb_instr_rt_idx_q_head_r_data = queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_instr_rt_idx__T_3_data = io_enq_0_bits_data_wb_instr_rt_idx;
  assign queue_bits_wb_instr_rt_idx__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_instr_rt_idx__T_3_mask = 1'h1;
  assign queue_bits_wb_instr_rt_idx__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_instr_rt_idx__T_4_data = io_enq_1_bits_data_wb_instr_rt_idx;
  assign queue_bits_wb_instr_rt_idx__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_instr_rt_idx__T_4_mask = 1'h1;
  assign queue_bits_wb_instr_rt_idx__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_instr_rt_idx__T_5_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_5_addr = 6'h0;
  assign queue_bits_wb_instr_rt_idx__T_5_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_5_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_6_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_6_addr = 6'h1;
  assign queue_bits_wb_instr_rt_idx__T_6_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_6_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_7_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_7_addr = 6'h2;
  assign queue_bits_wb_instr_rt_idx__T_7_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_7_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_8_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_8_addr = 6'h3;
  assign queue_bits_wb_instr_rt_idx__T_8_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_8_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_9_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_9_addr = 6'h4;
  assign queue_bits_wb_instr_rt_idx__T_9_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_9_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_10_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_10_addr = 6'h5;
  assign queue_bits_wb_instr_rt_idx__T_10_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_10_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_11_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_11_addr = 6'h6;
  assign queue_bits_wb_instr_rt_idx__T_11_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_11_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_12_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_12_addr = 6'h7;
  assign queue_bits_wb_instr_rt_idx__T_12_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_12_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_13_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_13_addr = 6'h8;
  assign queue_bits_wb_instr_rt_idx__T_13_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_13_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_14_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_14_addr = 6'h9;
  assign queue_bits_wb_instr_rt_idx__T_14_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_14_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_15_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_15_addr = 6'ha;
  assign queue_bits_wb_instr_rt_idx__T_15_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_15_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_16_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_16_addr = 6'hb;
  assign queue_bits_wb_instr_rt_idx__T_16_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_16_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_17_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_17_addr = 6'hc;
  assign queue_bits_wb_instr_rt_idx__T_17_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_17_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_18_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_18_addr = 6'hd;
  assign queue_bits_wb_instr_rt_idx__T_18_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_18_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_19_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_19_addr = 6'he;
  assign queue_bits_wb_instr_rt_idx__T_19_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_19_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_20_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_20_addr = 6'hf;
  assign queue_bits_wb_instr_rt_idx__T_20_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_20_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_21_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_21_addr = 6'h10;
  assign queue_bits_wb_instr_rt_idx__T_21_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_21_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_22_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_22_addr = 6'h11;
  assign queue_bits_wb_instr_rt_idx__T_22_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_22_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_23_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_23_addr = 6'h12;
  assign queue_bits_wb_instr_rt_idx__T_23_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_23_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_24_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_24_addr = 6'h13;
  assign queue_bits_wb_instr_rt_idx__T_24_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_24_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_25_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_25_addr = 6'h14;
  assign queue_bits_wb_instr_rt_idx__T_25_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_25_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_26_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_26_addr = 6'h15;
  assign queue_bits_wb_instr_rt_idx__T_26_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_26_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_27_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_27_addr = 6'h16;
  assign queue_bits_wb_instr_rt_idx__T_27_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_27_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_28_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_28_addr = 6'h17;
  assign queue_bits_wb_instr_rt_idx__T_28_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_28_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_29_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_29_addr = 6'h18;
  assign queue_bits_wb_instr_rt_idx__T_29_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_29_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_30_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_30_addr = 6'h19;
  assign queue_bits_wb_instr_rt_idx__T_30_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_30_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_31_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_31_addr = 6'h1a;
  assign queue_bits_wb_instr_rt_idx__T_31_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_31_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_32_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_32_addr = 6'h1b;
  assign queue_bits_wb_instr_rt_idx__T_32_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_32_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_33_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_33_addr = 6'h1c;
  assign queue_bits_wb_instr_rt_idx__T_33_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_33_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_34_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_34_addr = 6'h1d;
  assign queue_bits_wb_instr_rt_idx__T_34_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_34_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_35_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_35_addr = 6'h1e;
  assign queue_bits_wb_instr_rt_idx__T_35_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_35_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_36_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_36_addr = 6'h1f;
  assign queue_bits_wb_instr_rt_idx__T_36_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_36_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_37_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_37_addr = 6'h20;
  assign queue_bits_wb_instr_rt_idx__T_37_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_37_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_38_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_38_addr = 6'h21;
  assign queue_bits_wb_instr_rt_idx__T_38_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_38_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_39_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_39_addr = 6'h22;
  assign queue_bits_wb_instr_rt_idx__T_39_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_39_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_40_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_40_addr = 6'h23;
  assign queue_bits_wb_instr_rt_idx__T_40_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_40_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_41_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_41_addr = 6'h24;
  assign queue_bits_wb_instr_rt_idx__T_41_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_41_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_42_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_42_addr = 6'h25;
  assign queue_bits_wb_instr_rt_idx__T_42_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_42_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_43_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_43_addr = 6'h26;
  assign queue_bits_wb_instr_rt_idx__T_43_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_43_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_44_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_44_addr = 6'h27;
  assign queue_bits_wb_instr_rt_idx__T_44_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_44_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_45_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_45_addr = 6'h28;
  assign queue_bits_wb_instr_rt_idx__T_45_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_45_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_46_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_46_addr = 6'h29;
  assign queue_bits_wb_instr_rt_idx__T_46_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_46_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_47_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_47_addr = 6'h2a;
  assign queue_bits_wb_instr_rt_idx__T_47_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_47_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_48_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_48_addr = 6'h2b;
  assign queue_bits_wb_instr_rt_idx__T_48_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_48_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_49_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_49_addr = 6'h2c;
  assign queue_bits_wb_instr_rt_idx__T_49_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_49_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_50_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_50_addr = 6'h2d;
  assign queue_bits_wb_instr_rt_idx__T_50_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_50_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_51_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_51_addr = 6'h2e;
  assign queue_bits_wb_instr_rt_idx__T_51_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_51_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_52_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_52_addr = 6'h2f;
  assign queue_bits_wb_instr_rt_idx__T_52_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_52_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_53_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_53_addr = 6'h30;
  assign queue_bits_wb_instr_rt_idx__T_53_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_53_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_54_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_54_addr = 6'h31;
  assign queue_bits_wb_instr_rt_idx__T_54_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_54_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_55_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_55_addr = 6'h32;
  assign queue_bits_wb_instr_rt_idx__T_55_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_55_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_56_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_56_addr = 6'h33;
  assign queue_bits_wb_instr_rt_idx__T_56_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_56_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_57_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_57_addr = 6'h34;
  assign queue_bits_wb_instr_rt_idx__T_57_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_57_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_58_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_58_addr = 6'h35;
  assign queue_bits_wb_instr_rt_idx__T_58_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_58_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_59_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_59_addr = 6'h36;
  assign queue_bits_wb_instr_rt_idx__T_59_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_59_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_60_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_60_addr = 6'h37;
  assign queue_bits_wb_instr_rt_idx__T_60_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_60_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_61_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_61_addr = 6'h38;
  assign queue_bits_wb_instr_rt_idx__T_61_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_61_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_62_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_62_addr = 6'h39;
  assign queue_bits_wb_instr_rt_idx__T_62_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_62_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_63_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_63_addr = 6'h3a;
  assign queue_bits_wb_instr_rt_idx__T_63_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_63_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_64_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_64_addr = 6'h3b;
  assign queue_bits_wb_instr_rt_idx__T_64_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_64_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_65_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_65_addr = 6'h3c;
  assign queue_bits_wb_instr_rt_idx__T_65_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_65_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_66_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_66_addr = 6'h3d;
  assign queue_bits_wb_instr_rt_idx__T_66_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_66_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_67_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_67_addr = 6'h3e;
  assign queue_bits_wb_instr_rt_idx__T_67_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_67_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_68_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_68_addr = 6'h3f;
  assign queue_bits_wb_instr_rt_idx__T_68_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_68_en = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_70_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_70_addr = 6'h0;
  assign queue_bits_wb_instr_rt_idx__T_70_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_70_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_71_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_71_addr = 6'h1;
  assign queue_bits_wb_instr_rt_idx__T_71_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_71_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_72_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_72_addr = 6'h2;
  assign queue_bits_wb_instr_rt_idx__T_72_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_72_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_73_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_73_addr = 6'h3;
  assign queue_bits_wb_instr_rt_idx__T_73_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_73_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_74_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_74_addr = 6'h4;
  assign queue_bits_wb_instr_rt_idx__T_74_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_74_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_75_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_75_addr = 6'h5;
  assign queue_bits_wb_instr_rt_idx__T_75_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_75_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_76_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_76_addr = 6'h6;
  assign queue_bits_wb_instr_rt_idx__T_76_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_76_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_77_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_77_addr = 6'h7;
  assign queue_bits_wb_instr_rt_idx__T_77_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_77_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_78_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_78_addr = 6'h8;
  assign queue_bits_wb_instr_rt_idx__T_78_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_78_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_79_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_79_addr = 6'h9;
  assign queue_bits_wb_instr_rt_idx__T_79_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_79_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_80_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_80_addr = 6'ha;
  assign queue_bits_wb_instr_rt_idx__T_80_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_80_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_81_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_81_addr = 6'hb;
  assign queue_bits_wb_instr_rt_idx__T_81_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_81_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_82_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_82_addr = 6'hc;
  assign queue_bits_wb_instr_rt_idx__T_82_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_82_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_83_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_83_addr = 6'hd;
  assign queue_bits_wb_instr_rt_idx__T_83_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_83_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_84_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_84_addr = 6'he;
  assign queue_bits_wb_instr_rt_idx__T_84_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_84_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_85_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_85_addr = 6'hf;
  assign queue_bits_wb_instr_rt_idx__T_85_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_85_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_86_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_86_addr = 6'h10;
  assign queue_bits_wb_instr_rt_idx__T_86_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_86_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_87_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_87_addr = 6'h11;
  assign queue_bits_wb_instr_rt_idx__T_87_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_87_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_88_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_88_addr = 6'h12;
  assign queue_bits_wb_instr_rt_idx__T_88_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_88_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_89_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_89_addr = 6'h13;
  assign queue_bits_wb_instr_rt_idx__T_89_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_89_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_90_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_90_addr = 6'h14;
  assign queue_bits_wb_instr_rt_idx__T_90_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_90_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_91_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_91_addr = 6'h15;
  assign queue_bits_wb_instr_rt_idx__T_91_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_91_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_92_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_92_addr = 6'h16;
  assign queue_bits_wb_instr_rt_idx__T_92_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_92_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_93_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_93_addr = 6'h17;
  assign queue_bits_wb_instr_rt_idx__T_93_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_93_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_94_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_94_addr = 6'h18;
  assign queue_bits_wb_instr_rt_idx__T_94_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_94_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_95_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_95_addr = 6'h19;
  assign queue_bits_wb_instr_rt_idx__T_95_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_95_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_96_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_96_addr = 6'h1a;
  assign queue_bits_wb_instr_rt_idx__T_96_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_96_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_97_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_97_addr = 6'h1b;
  assign queue_bits_wb_instr_rt_idx__T_97_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_97_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_98_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_98_addr = 6'h1c;
  assign queue_bits_wb_instr_rt_idx__T_98_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_98_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_99_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_99_addr = 6'h1d;
  assign queue_bits_wb_instr_rt_idx__T_99_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_99_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_100_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_100_addr = 6'h1e;
  assign queue_bits_wb_instr_rt_idx__T_100_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_100_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_101_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_101_addr = 6'h1f;
  assign queue_bits_wb_instr_rt_idx__T_101_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_101_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_102_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_102_addr = 6'h20;
  assign queue_bits_wb_instr_rt_idx__T_102_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_102_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_103_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_103_addr = 6'h21;
  assign queue_bits_wb_instr_rt_idx__T_103_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_103_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_104_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_104_addr = 6'h22;
  assign queue_bits_wb_instr_rt_idx__T_104_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_104_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_105_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_105_addr = 6'h23;
  assign queue_bits_wb_instr_rt_idx__T_105_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_105_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_106_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_106_addr = 6'h24;
  assign queue_bits_wb_instr_rt_idx__T_106_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_106_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_107_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_107_addr = 6'h25;
  assign queue_bits_wb_instr_rt_idx__T_107_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_107_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_108_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_108_addr = 6'h26;
  assign queue_bits_wb_instr_rt_idx__T_108_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_108_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_109_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_109_addr = 6'h27;
  assign queue_bits_wb_instr_rt_idx__T_109_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_109_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_110_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_110_addr = 6'h28;
  assign queue_bits_wb_instr_rt_idx__T_110_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_110_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_111_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_111_addr = 6'h29;
  assign queue_bits_wb_instr_rt_idx__T_111_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_111_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_112_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_112_addr = 6'h2a;
  assign queue_bits_wb_instr_rt_idx__T_112_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_112_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_113_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_113_addr = 6'h2b;
  assign queue_bits_wb_instr_rt_idx__T_113_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_113_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_114_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_114_addr = 6'h2c;
  assign queue_bits_wb_instr_rt_idx__T_114_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_114_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_115_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_115_addr = 6'h2d;
  assign queue_bits_wb_instr_rt_idx__T_115_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_115_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_116_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_116_addr = 6'h2e;
  assign queue_bits_wb_instr_rt_idx__T_116_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_116_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_117_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_117_addr = 6'h2f;
  assign queue_bits_wb_instr_rt_idx__T_117_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_117_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_118_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_118_addr = 6'h30;
  assign queue_bits_wb_instr_rt_idx__T_118_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_118_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_119_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_119_addr = 6'h31;
  assign queue_bits_wb_instr_rt_idx__T_119_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_119_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_120_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_120_addr = 6'h32;
  assign queue_bits_wb_instr_rt_idx__T_120_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_120_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_121_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_121_addr = 6'h33;
  assign queue_bits_wb_instr_rt_idx__T_121_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_121_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_122_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_122_addr = 6'h34;
  assign queue_bits_wb_instr_rt_idx__T_122_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_122_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_123_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_123_addr = 6'h35;
  assign queue_bits_wb_instr_rt_idx__T_123_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_123_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_124_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_124_addr = 6'h36;
  assign queue_bits_wb_instr_rt_idx__T_124_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_124_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_125_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_125_addr = 6'h37;
  assign queue_bits_wb_instr_rt_idx__T_125_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_125_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_126_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_126_addr = 6'h38;
  assign queue_bits_wb_instr_rt_idx__T_126_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_126_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_127_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_127_addr = 6'h39;
  assign queue_bits_wb_instr_rt_idx__T_127_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_127_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_128_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_128_addr = 6'h3a;
  assign queue_bits_wb_instr_rt_idx__T_128_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_128_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_129_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_129_addr = 6'h3b;
  assign queue_bits_wb_instr_rt_idx__T_129_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_129_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_130_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_130_addr = 6'h3c;
  assign queue_bits_wb_instr_rt_idx__T_130_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_130_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_131_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_131_addr = 6'h3d;
  assign queue_bits_wb_instr_rt_idx__T_131_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_131_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_132_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_132_addr = 6'h3e;
  assign queue_bits_wb_instr_rt_idx__T_132_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_132_en = reset;
  assign queue_bits_wb_instr_rt_idx__T_133_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx__T_133_addr = 6'h3f;
  assign queue_bits_wb_instr_rt_idx__T_133_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx__T_133_en = reset;
  assign queue_bits_wb_instr_rt_idx_q_head_w_data = 5'h0;
  assign queue_bits_wb_instr_rt_idx_q_head_w_addr = head;
  assign queue_bits_wb_instr_rt_idx_q_head_w_mask = 1'h0;
  assign queue_bits_wb_instr_rt_idx_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_instr_rd_idx_q_head_r_addr = head;
  assign queue_bits_wb_instr_rd_idx_q_head_r_data = queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_instr_rd_idx__T_3_data = io_enq_0_bits_data_wb_instr_rd_idx;
  assign queue_bits_wb_instr_rd_idx__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_instr_rd_idx__T_3_mask = 1'h1;
  assign queue_bits_wb_instr_rd_idx__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_instr_rd_idx__T_4_data = io_enq_1_bits_data_wb_instr_rd_idx;
  assign queue_bits_wb_instr_rd_idx__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_instr_rd_idx__T_4_mask = 1'h1;
  assign queue_bits_wb_instr_rd_idx__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_instr_rd_idx__T_5_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_5_addr = 6'h0;
  assign queue_bits_wb_instr_rd_idx__T_5_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_5_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_6_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_6_addr = 6'h1;
  assign queue_bits_wb_instr_rd_idx__T_6_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_6_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_7_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_7_addr = 6'h2;
  assign queue_bits_wb_instr_rd_idx__T_7_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_7_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_8_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_8_addr = 6'h3;
  assign queue_bits_wb_instr_rd_idx__T_8_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_8_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_9_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_9_addr = 6'h4;
  assign queue_bits_wb_instr_rd_idx__T_9_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_9_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_10_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_10_addr = 6'h5;
  assign queue_bits_wb_instr_rd_idx__T_10_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_10_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_11_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_11_addr = 6'h6;
  assign queue_bits_wb_instr_rd_idx__T_11_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_11_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_12_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_12_addr = 6'h7;
  assign queue_bits_wb_instr_rd_idx__T_12_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_12_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_13_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_13_addr = 6'h8;
  assign queue_bits_wb_instr_rd_idx__T_13_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_13_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_14_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_14_addr = 6'h9;
  assign queue_bits_wb_instr_rd_idx__T_14_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_14_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_15_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_15_addr = 6'ha;
  assign queue_bits_wb_instr_rd_idx__T_15_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_15_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_16_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_16_addr = 6'hb;
  assign queue_bits_wb_instr_rd_idx__T_16_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_16_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_17_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_17_addr = 6'hc;
  assign queue_bits_wb_instr_rd_idx__T_17_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_17_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_18_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_18_addr = 6'hd;
  assign queue_bits_wb_instr_rd_idx__T_18_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_18_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_19_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_19_addr = 6'he;
  assign queue_bits_wb_instr_rd_idx__T_19_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_19_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_20_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_20_addr = 6'hf;
  assign queue_bits_wb_instr_rd_idx__T_20_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_20_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_21_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_21_addr = 6'h10;
  assign queue_bits_wb_instr_rd_idx__T_21_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_21_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_22_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_22_addr = 6'h11;
  assign queue_bits_wb_instr_rd_idx__T_22_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_22_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_23_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_23_addr = 6'h12;
  assign queue_bits_wb_instr_rd_idx__T_23_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_23_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_24_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_24_addr = 6'h13;
  assign queue_bits_wb_instr_rd_idx__T_24_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_24_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_25_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_25_addr = 6'h14;
  assign queue_bits_wb_instr_rd_idx__T_25_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_25_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_26_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_26_addr = 6'h15;
  assign queue_bits_wb_instr_rd_idx__T_26_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_26_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_27_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_27_addr = 6'h16;
  assign queue_bits_wb_instr_rd_idx__T_27_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_27_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_28_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_28_addr = 6'h17;
  assign queue_bits_wb_instr_rd_idx__T_28_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_28_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_29_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_29_addr = 6'h18;
  assign queue_bits_wb_instr_rd_idx__T_29_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_29_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_30_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_30_addr = 6'h19;
  assign queue_bits_wb_instr_rd_idx__T_30_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_30_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_31_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_31_addr = 6'h1a;
  assign queue_bits_wb_instr_rd_idx__T_31_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_31_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_32_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_32_addr = 6'h1b;
  assign queue_bits_wb_instr_rd_idx__T_32_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_32_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_33_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_33_addr = 6'h1c;
  assign queue_bits_wb_instr_rd_idx__T_33_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_33_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_34_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_34_addr = 6'h1d;
  assign queue_bits_wb_instr_rd_idx__T_34_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_34_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_35_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_35_addr = 6'h1e;
  assign queue_bits_wb_instr_rd_idx__T_35_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_35_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_36_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_36_addr = 6'h1f;
  assign queue_bits_wb_instr_rd_idx__T_36_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_36_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_37_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_37_addr = 6'h20;
  assign queue_bits_wb_instr_rd_idx__T_37_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_37_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_38_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_38_addr = 6'h21;
  assign queue_bits_wb_instr_rd_idx__T_38_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_38_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_39_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_39_addr = 6'h22;
  assign queue_bits_wb_instr_rd_idx__T_39_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_39_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_40_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_40_addr = 6'h23;
  assign queue_bits_wb_instr_rd_idx__T_40_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_40_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_41_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_41_addr = 6'h24;
  assign queue_bits_wb_instr_rd_idx__T_41_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_41_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_42_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_42_addr = 6'h25;
  assign queue_bits_wb_instr_rd_idx__T_42_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_42_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_43_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_43_addr = 6'h26;
  assign queue_bits_wb_instr_rd_idx__T_43_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_43_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_44_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_44_addr = 6'h27;
  assign queue_bits_wb_instr_rd_idx__T_44_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_44_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_45_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_45_addr = 6'h28;
  assign queue_bits_wb_instr_rd_idx__T_45_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_45_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_46_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_46_addr = 6'h29;
  assign queue_bits_wb_instr_rd_idx__T_46_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_46_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_47_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_47_addr = 6'h2a;
  assign queue_bits_wb_instr_rd_idx__T_47_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_47_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_48_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_48_addr = 6'h2b;
  assign queue_bits_wb_instr_rd_idx__T_48_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_48_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_49_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_49_addr = 6'h2c;
  assign queue_bits_wb_instr_rd_idx__T_49_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_49_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_50_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_50_addr = 6'h2d;
  assign queue_bits_wb_instr_rd_idx__T_50_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_50_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_51_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_51_addr = 6'h2e;
  assign queue_bits_wb_instr_rd_idx__T_51_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_51_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_52_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_52_addr = 6'h2f;
  assign queue_bits_wb_instr_rd_idx__T_52_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_52_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_53_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_53_addr = 6'h30;
  assign queue_bits_wb_instr_rd_idx__T_53_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_53_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_54_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_54_addr = 6'h31;
  assign queue_bits_wb_instr_rd_idx__T_54_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_54_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_55_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_55_addr = 6'h32;
  assign queue_bits_wb_instr_rd_idx__T_55_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_55_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_56_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_56_addr = 6'h33;
  assign queue_bits_wb_instr_rd_idx__T_56_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_56_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_57_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_57_addr = 6'h34;
  assign queue_bits_wb_instr_rd_idx__T_57_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_57_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_58_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_58_addr = 6'h35;
  assign queue_bits_wb_instr_rd_idx__T_58_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_58_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_59_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_59_addr = 6'h36;
  assign queue_bits_wb_instr_rd_idx__T_59_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_59_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_60_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_60_addr = 6'h37;
  assign queue_bits_wb_instr_rd_idx__T_60_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_60_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_61_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_61_addr = 6'h38;
  assign queue_bits_wb_instr_rd_idx__T_61_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_61_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_62_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_62_addr = 6'h39;
  assign queue_bits_wb_instr_rd_idx__T_62_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_62_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_63_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_63_addr = 6'h3a;
  assign queue_bits_wb_instr_rd_idx__T_63_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_63_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_64_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_64_addr = 6'h3b;
  assign queue_bits_wb_instr_rd_idx__T_64_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_64_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_65_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_65_addr = 6'h3c;
  assign queue_bits_wb_instr_rd_idx__T_65_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_65_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_66_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_66_addr = 6'h3d;
  assign queue_bits_wb_instr_rd_idx__T_66_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_66_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_67_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_67_addr = 6'h3e;
  assign queue_bits_wb_instr_rd_idx__T_67_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_67_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_68_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_68_addr = 6'h3f;
  assign queue_bits_wb_instr_rd_idx__T_68_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_68_en = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_70_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_70_addr = 6'h0;
  assign queue_bits_wb_instr_rd_idx__T_70_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_70_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_71_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_71_addr = 6'h1;
  assign queue_bits_wb_instr_rd_idx__T_71_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_71_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_72_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_72_addr = 6'h2;
  assign queue_bits_wb_instr_rd_idx__T_72_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_72_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_73_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_73_addr = 6'h3;
  assign queue_bits_wb_instr_rd_idx__T_73_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_73_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_74_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_74_addr = 6'h4;
  assign queue_bits_wb_instr_rd_idx__T_74_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_74_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_75_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_75_addr = 6'h5;
  assign queue_bits_wb_instr_rd_idx__T_75_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_75_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_76_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_76_addr = 6'h6;
  assign queue_bits_wb_instr_rd_idx__T_76_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_76_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_77_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_77_addr = 6'h7;
  assign queue_bits_wb_instr_rd_idx__T_77_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_77_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_78_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_78_addr = 6'h8;
  assign queue_bits_wb_instr_rd_idx__T_78_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_78_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_79_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_79_addr = 6'h9;
  assign queue_bits_wb_instr_rd_idx__T_79_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_79_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_80_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_80_addr = 6'ha;
  assign queue_bits_wb_instr_rd_idx__T_80_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_80_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_81_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_81_addr = 6'hb;
  assign queue_bits_wb_instr_rd_idx__T_81_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_81_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_82_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_82_addr = 6'hc;
  assign queue_bits_wb_instr_rd_idx__T_82_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_82_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_83_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_83_addr = 6'hd;
  assign queue_bits_wb_instr_rd_idx__T_83_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_83_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_84_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_84_addr = 6'he;
  assign queue_bits_wb_instr_rd_idx__T_84_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_84_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_85_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_85_addr = 6'hf;
  assign queue_bits_wb_instr_rd_idx__T_85_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_85_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_86_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_86_addr = 6'h10;
  assign queue_bits_wb_instr_rd_idx__T_86_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_86_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_87_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_87_addr = 6'h11;
  assign queue_bits_wb_instr_rd_idx__T_87_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_87_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_88_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_88_addr = 6'h12;
  assign queue_bits_wb_instr_rd_idx__T_88_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_88_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_89_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_89_addr = 6'h13;
  assign queue_bits_wb_instr_rd_idx__T_89_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_89_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_90_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_90_addr = 6'h14;
  assign queue_bits_wb_instr_rd_idx__T_90_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_90_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_91_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_91_addr = 6'h15;
  assign queue_bits_wb_instr_rd_idx__T_91_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_91_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_92_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_92_addr = 6'h16;
  assign queue_bits_wb_instr_rd_idx__T_92_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_92_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_93_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_93_addr = 6'h17;
  assign queue_bits_wb_instr_rd_idx__T_93_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_93_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_94_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_94_addr = 6'h18;
  assign queue_bits_wb_instr_rd_idx__T_94_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_94_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_95_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_95_addr = 6'h19;
  assign queue_bits_wb_instr_rd_idx__T_95_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_95_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_96_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_96_addr = 6'h1a;
  assign queue_bits_wb_instr_rd_idx__T_96_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_96_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_97_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_97_addr = 6'h1b;
  assign queue_bits_wb_instr_rd_idx__T_97_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_97_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_98_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_98_addr = 6'h1c;
  assign queue_bits_wb_instr_rd_idx__T_98_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_98_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_99_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_99_addr = 6'h1d;
  assign queue_bits_wb_instr_rd_idx__T_99_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_99_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_100_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_100_addr = 6'h1e;
  assign queue_bits_wb_instr_rd_idx__T_100_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_100_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_101_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_101_addr = 6'h1f;
  assign queue_bits_wb_instr_rd_idx__T_101_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_101_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_102_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_102_addr = 6'h20;
  assign queue_bits_wb_instr_rd_idx__T_102_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_102_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_103_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_103_addr = 6'h21;
  assign queue_bits_wb_instr_rd_idx__T_103_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_103_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_104_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_104_addr = 6'h22;
  assign queue_bits_wb_instr_rd_idx__T_104_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_104_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_105_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_105_addr = 6'h23;
  assign queue_bits_wb_instr_rd_idx__T_105_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_105_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_106_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_106_addr = 6'h24;
  assign queue_bits_wb_instr_rd_idx__T_106_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_106_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_107_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_107_addr = 6'h25;
  assign queue_bits_wb_instr_rd_idx__T_107_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_107_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_108_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_108_addr = 6'h26;
  assign queue_bits_wb_instr_rd_idx__T_108_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_108_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_109_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_109_addr = 6'h27;
  assign queue_bits_wb_instr_rd_idx__T_109_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_109_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_110_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_110_addr = 6'h28;
  assign queue_bits_wb_instr_rd_idx__T_110_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_110_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_111_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_111_addr = 6'h29;
  assign queue_bits_wb_instr_rd_idx__T_111_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_111_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_112_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_112_addr = 6'h2a;
  assign queue_bits_wb_instr_rd_idx__T_112_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_112_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_113_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_113_addr = 6'h2b;
  assign queue_bits_wb_instr_rd_idx__T_113_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_113_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_114_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_114_addr = 6'h2c;
  assign queue_bits_wb_instr_rd_idx__T_114_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_114_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_115_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_115_addr = 6'h2d;
  assign queue_bits_wb_instr_rd_idx__T_115_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_115_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_116_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_116_addr = 6'h2e;
  assign queue_bits_wb_instr_rd_idx__T_116_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_116_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_117_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_117_addr = 6'h2f;
  assign queue_bits_wb_instr_rd_idx__T_117_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_117_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_118_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_118_addr = 6'h30;
  assign queue_bits_wb_instr_rd_idx__T_118_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_118_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_119_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_119_addr = 6'h31;
  assign queue_bits_wb_instr_rd_idx__T_119_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_119_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_120_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_120_addr = 6'h32;
  assign queue_bits_wb_instr_rd_idx__T_120_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_120_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_121_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_121_addr = 6'h33;
  assign queue_bits_wb_instr_rd_idx__T_121_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_121_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_122_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_122_addr = 6'h34;
  assign queue_bits_wb_instr_rd_idx__T_122_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_122_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_123_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_123_addr = 6'h35;
  assign queue_bits_wb_instr_rd_idx__T_123_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_123_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_124_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_124_addr = 6'h36;
  assign queue_bits_wb_instr_rd_idx__T_124_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_124_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_125_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_125_addr = 6'h37;
  assign queue_bits_wb_instr_rd_idx__T_125_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_125_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_126_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_126_addr = 6'h38;
  assign queue_bits_wb_instr_rd_idx__T_126_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_126_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_127_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_127_addr = 6'h39;
  assign queue_bits_wb_instr_rd_idx__T_127_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_127_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_128_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_128_addr = 6'h3a;
  assign queue_bits_wb_instr_rd_idx__T_128_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_128_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_129_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_129_addr = 6'h3b;
  assign queue_bits_wb_instr_rd_idx__T_129_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_129_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_130_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_130_addr = 6'h3c;
  assign queue_bits_wb_instr_rd_idx__T_130_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_130_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_131_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_131_addr = 6'h3d;
  assign queue_bits_wb_instr_rd_idx__T_131_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_131_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_132_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_132_addr = 6'h3e;
  assign queue_bits_wb_instr_rd_idx__T_132_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_132_en = reset;
  assign queue_bits_wb_instr_rd_idx__T_133_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx__T_133_addr = 6'h3f;
  assign queue_bits_wb_instr_rd_idx__T_133_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx__T_133_en = reset;
  assign queue_bits_wb_instr_rd_idx_q_head_w_data = 5'h0;
  assign queue_bits_wb_instr_rd_idx_q_head_w_addr = head;
  assign queue_bits_wb_instr_rd_idx_q_head_w_mask = 1'h0;
  assign queue_bits_wb_instr_rd_idx_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_instr_shamt_q_head_r_addr = head;
  assign queue_bits_wb_instr_shamt_q_head_r_data = queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_instr_shamt__T_3_data = io_enq_0_bits_data_wb_instr_shamt;
  assign queue_bits_wb_instr_shamt__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_instr_shamt__T_3_mask = 1'h1;
  assign queue_bits_wb_instr_shamt__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_instr_shamt__T_4_data = io_enq_1_bits_data_wb_instr_shamt;
  assign queue_bits_wb_instr_shamt__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_instr_shamt__T_4_mask = 1'h1;
  assign queue_bits_wb_instr_shamt__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_instr_shamt__T_5_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_5_addr = 6'h0;
  assign queue_bits_wb_instr_shamt__T_5_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_5_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_6_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_6_addr = 6'h1;
  assign queue_bits_wb_instr_shamt__T_6_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_6_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_7_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_7_addr = 6'h2;
  assign queue_bits_wb_instr_shamt__T_7_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_7_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_8_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_8_addr = 6'h3;
  assign queue_bits_wb_instr_shamt__T_8_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_8_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_9_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_9_addr = 6'h4;
  assign queue_bits_wb_instr_shamt__T_9_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_9_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_10_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_10_addr = 6'h5;
  assign queue_bits_wb_instr_shamt__T_10_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_10_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_11_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_11_addr = 6'h6;
  assign queue_bits_wb_instr_shamt__T_11_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_11_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_12_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_12_addr = 6'h7;
  assign queue_bits_wb_instr_shamt__T_12_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_12_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_13_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_13_addr = 6'h8;
  assign queue_bits_wb_instr_shamt__T_13_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_13_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_14_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_14_addr = 6'h9;
  assign queue_bits_wb_instr_shamt__T_14_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_14_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_15_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_15_addr = 6'ha;
  assign queue_bits_wb_instr_shamt__T_15_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_15_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_16_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_16_addr = 6'hb;
  assign queue_bits_wb_instr_shamt__T_16_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_16_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_17_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_17_addr = 6'hc;
  assign queue_bits_wb_instr_shamt__T_17_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_17_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_18_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_18_addr = 6'hd;
  assign queue_bits_wb_instr_shamt__T_18_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_18_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_19_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_19_addr = 6'he;
  assign queue_bits_wb_instr_shamt__T_19_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_19_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_20_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_20_addr = 6'hf;
  assign queue_bits_wb_instr_shamt__T_20_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_20_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_21_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_21_addr = 6'h10;
  assign queue_bits_wb_instr_shamt__T_21_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_21_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_22_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_22_addr = 6'h11;
  assign queue_bits_wb_instr_shamt__T_22_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_22_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_23_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_23_addr = 6'h12;
  assign queue_bits_wb_instr_shamt__T_23_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_23_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_24_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_24_addr = 6'h13;
  assign queue_bits_wb_instr_shamt__T_24_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_24_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_25_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_25_addr = 6'h14;
  assign queue_bits_wb_instr_shamt__T_25_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_25_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_26_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_26_addr = 6'h15;
  assign queue_bits_wb_instr_shamt__T_26_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_26_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_27_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_27_addr = 6'h16;
  assign queue_bits_wb_instr_shamt__T_27_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_27_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_28_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_28_addr = 6'h17;
  assign queue_bits_wb_instr_shamt__T_28_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_28_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_29_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_29_addr = 6'h18;
  assign queue_bits_wb_instr_shamt__T_29_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_29_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_30_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_30_addr = 6'h19;
  assign queue_bits_wb_instr_shamt__T_30_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_30_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_31_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_31_addr = 6'h1a;
  assign queue_bits_wb_instr_shamt__T_31_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_31_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_32_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_32_addr = 6'h1b;
  assign queue_bits_wb_instr_shamt__T_32_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_32_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_33_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_33_addr = 6'h1c;
  assign queue_bits_wb_instr_shamt__T_33_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_33_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_34_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_34_addr = 6'h1d;
  assign queue_bits_wb_instr_shamt__T_34_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_34_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_35_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_35_addr = 6'h1e;
  assign queue_bits_wb_instr_shamt__T_35_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_35_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_36_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_36_addr = 6'h1f;
  assign queue_bits_wb_instr_shamt__T_36_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_36_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_37_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_37_addr = 6'h20;
  assign queue_bits_wb_instr_shamt__T_37_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_37_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_38_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_38_addr = 6'h21;
  assign queue_bits_wb_instr_shamt__T_38_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_38_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_39_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_39_addr = 6'h22;
  assign queue_bits_wb_instr_shamt__T_39_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_39_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_40_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_40_addr = 6'h23;
  assign queue_bits_wb_instr_shamt__T_40_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_40_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_41_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_41_addr = 6'h24;
  assign queue_bits_wb_instr_shamt__T_41_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_41_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_42_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_42_addr = 6'h25;
  assign queue_bits_wb_instr_shamt__T_42_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_42_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_43_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_43_addr = 6'h26;
  assign queue_bits_wb_instr_shamt__T_43_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_43_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_44_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_44_addr = 6'h27;
  assign queue_bits_wb_instr_shamt__T_44_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_44_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_45_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_45_addr = 6'h28;
  assign queue_bits_wb_instr_shamt__T_45_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_45_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_46_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_46_addr = 6'h29;
  assign queue_bits_wb_instr_shamt__T_46_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_46_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_47_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_47_addr = 6'h2a;
  assign queue_bits_wb_instr_shamt__T_47_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_47_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_48_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_48_addr = 6'h2b;
  assign queue_bits_wb_instr_shamt__T_48_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_48_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_49_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_49_addr = 6'h2c;
  assign queue_bits_wb_instr_shamt__T_49_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_49_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_50_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_50_addr = 6'h2d;
  assign queue_bits_wb_instr_shamt__T_50_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_50_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_51_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_51_addr = 6'h2e;
  assign queue_bits_wb_instr_shamt__T_51_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_51_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_52_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_52_addr = 6'h2f;
  assign queue_bits_wb_instr_shamt__T_52_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_52_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_53_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_53_addr = 6'h30;
  assign queue_bits_wb_instr_shamt__T_53_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_53_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_54_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_54_addr = 6'h31;
  assign queue_bits_wb_instr_shamt__T_54_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_54_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_55_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_55_addr = 6'h32;
  assign queue_bits_wb_instr_shamt__T_55_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_55_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_56_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_56_addr = 6'h33;
  assign queue_bits_wb_instr_shamt__T_56_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_56_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_57_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_57_addr = 6'h34;
  assign queue_bits_wb_instr_shamt__T_57_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_57_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_58_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_58_addr = 6'h35;
  assign queue_bits_wb_instr_shamt__T_58_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_58_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_59_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_59_addr = 6'h36;
  assign queue_bits_wb_instr_shamt__T_59_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_59_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_60_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_60_addr = 6'h37;
  assign queue_bits_wb_instr_shamt__T_60_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_60_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_61_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_61_addr = 6'h38;
  assign queue_bits_wb_instr_shamt__T_61_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_61_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_62_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_62_addr = 6'h39;
  assign queue_bits_wb_instr_shamt__T_62_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_62_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_63_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_63_addr = 6'h3a;
  assign queue_bits_wb_instr_shamt__T_63_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_63_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_64_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_64_addr = 6'h3b;
  assign queue_bits_wb_instr_shamt__T_64_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_64_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_65_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_65_addr = 6'h3c;
  assign queue_bits_wb_instr_shamt__T_65_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_65_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_66_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_66_addr = 6'h3d;
  assign queue_bits_wb_instr_shamt__T_66_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_66_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_67_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_67_addr = 6'h3e;
  assign queue_bits_wb_instr_shamt__T_67_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_67_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_68_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_68_addr = 6'h3f;
  assign queue_bits_wb_instr_shamt__T_68_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_68_en = 1'h0;
  assign queue_bits_wb_instr_shamt__T_70_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_70_addr = 6'h0;
  assign queue_bits_wb_instr_shamt__T_70_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_70_en = reset;
  assign queue_bits_wb_instr_shamt__T_71_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_71_addr = 6'h1;
  assign queue_bits_wb_instr_shamt__T_71_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_71_en = reset;
  assign queue_bits_wb_instr_shamt__T_72_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_72_addr = 6'h2;
  assign queue_bits_wb_instr_shamt__T_72_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_72_en = reset;
  assign queue_bits_wb_instr_shamt__T_73_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_73_addr = 6'h3;
  assign queue_bits_wb_instr_shamt__T_73_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_73_en = reset;
  assign queue_bits_wb_instr_shamt__T_74_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_74_addr = 6'h4;
  assign queue_bits_wb_instr_shamt__T_74_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_74_en = reset;
  assign queue_bits_wb_instr_shamt__T_75_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_75_addr = 6'h5;
  assign queue_bits_wb_instr_shamt__T_75_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_75_en = reset;
  assign queue_bits_wb_instr_shamt__T_76_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_76_addr = 6'h6;
  assign queue_bits_wb_instr_shamt__T_76_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_76_en = reset;
  assign queue_bits_wb_instr_shamt__T_77_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_77_addr = 6'h7;
  assign queue_bits_wb_instr_shamt__T_77_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_77_en = reset;
  assign queue_bits_wb_instr_shamt__T_78_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_78_addr = 6'h8;
  assign queue_bits_wb_instr_shamt__T_78_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_78_en = reset;
  assign queue_bits_wb_instr_shamt__T_79_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_79_addr = 6'h9;
  assign queue_bits_wb_instr_shamt__T_79_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_79_en = reset;
  assign queue_bits_wb_instr_shamt__T_80_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_80_addr = 6'ha;
  assign queue_bits_wb_instr_shamt__T_80_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_80_en = reset;
  assign queue_bits_wb_instr_shamt__T_81_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_81_addr = 6'hb;
  assign queue_bits_wb_instr_shamt__T_81_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_81_en = reset;
  assign queue_bits_wb_instr_shamt__T_82_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_82_addr = 6'hc;
  assign queue_bits_wb_instr_shamt__T_82_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_82_en = reset;
  assign queue_bits_wb_instr_shamt__T_83_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_83_addr = 6'hd;
  assign queue_bits_wb_instr_shamt__T_83_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_83_en = reset;
  assign queue_bits_wb_instr_shamt__T_84_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_84_addr = 6'he;
  assign queue_bits_wb_instr_shamt__T_84_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_84_en = reset;
  assign queue_bits_wb_instr_shamt__T_85_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_85_addr = 6'hf;
  assign queue_bits_wb_instr_shamt__T_85_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_85_en = reset;
  assign queue_bits_wb_instr_shamt__T_86_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_86_addr = 6'h10;
  assign queue_bits_wb_instr_shamt__T_86_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_86_en = reset;
  assign queue_bits_wb_instr_shamt__T_87_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_87_addr = 6'h11;
  assign queue_bits_wb_instr_shamt__T_87_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_87_en = reset;
  assign queue_bits_wb_instr_shamt__T_88_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_88_addr = 6'h12;
  assign queue_bits_wb_instr_shamt__T_88_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_88_en = reset;
  assign queue_bits_wb_instr_shamt__T_89_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_89_addr = 6'h13;
  assign queue_bits_wb_instr_shamt__T_89_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_89_en = reset;
  assign queue_bits_wb_instr_shamt__T_90_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_90_addr = 6'h14;
  assign queue_bits_wb_instr_shamt__T_90_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_90_en = reset;
  assign queue_bits_wb_instr_shamt__T_91_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_91_addr = 6'h15;
  assign queue_bits_wb_instr_shamt__T_91_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_91_en = reset;
  assign queue_bits_wb_instr_shamt__T_92_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_92_addr = 6'h16;
  assign queue_bits_wb_instr_shamt__T_92_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_92_en = reset;
  assign queue_bits_wb_instr_shamt__T_93_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_93_addr = 6'h17;
  assign queue_bits_wb_instr_shamt__T_93_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_93_en = reset;
  assign queue_bits_wb_instr_shamt__T_94_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_94_addr = 6'h18;
  assign queue_bits_wb_instr_shamt__T_94_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_94_en = reset;
  assign queue_bits_wb_instr_shamt__T_95_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_95_addr = 6'h19;
  assign queue_bits_wb_instr_shamt__T_95_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_95_en = reset;
  assign queue_bits_wb_instr_shamt__T_96_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_96_addr = 6'h1a;
  assign queue_bits_wb_instr_shamt__T_96_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_96_en = reset;
  assign queue_bits_wb_instr_shamt__T_97_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_97_addr = 6'h1b;
  assign queue_bits_wb_instr_shamt__T_97_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_97_en = reset;
  assign queue_bits_wb_instr_shamt__T_98_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_98_addr = 6'h1c;
  assign queue_bits_wb_instr_shamt__T_98_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_98_en = reset;
  assign queue_bits_wb_instr_shamt__T_99_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_99_addr = 6'h1d;
  assign queue_bits_wb_instr_shamt__T_99_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_99_en = reset;
  assign queue_bits_wb_instr_shamt__T_100_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_100_addr = 6'h1e;
  assign queue_bits_wb_instr_shamt__T_100_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_100_en = reset;
  assign queue_bits_wb_instr_shamt__T_101_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_101_addr = 6'h1f;
  assign queue_bits_wb_instr_shamt__T_101_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_101_en = reset;
  assign queue_bits_wb_instr_shamt__T_102_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_102_addr = 6'h20;
  assign queue_bits_wb_instr_shamt__T_102_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_102_en = reset;
  assign queue_bits_wb_instr_shamt__T_103_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_103_addr = 6'h21;
  assign queue_bits_wb_instr_shamt__T_103_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_103_en = reset;
  assign queue_bits_wb_instr_shamt__T_104_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_104_addr = 6'h22;
  assign queue_bits_wb_instr_shamt__T_104_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_104_en = reset;
  assign queue_bits_wb_instr_shamt__T_105_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_105_addr = 6'h23;
  assign queue_bits_wb_instr_shamt__T_105_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_105_en = reset;
  assign queue_bits_wb_instr_shamt__T_106_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_106_addr = 6'h24;
  assign queue_bits_wb_instr_shamt__T_106_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_106_en = reset;
  assign queue_bits_wb_instr_shamt__T_107_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_107_addr = 6'h25;
  assign queue_bits_wb_instr_shamt__T_107_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_107_en = reset;
  assign queue_bits_wb_instr_shamt__T_108_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_108_addr = 6'h26;
  assign queue_bits_wb_instr_shamt__T_108_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_108_en = reset;
  assign queue_bits_wb_instr_shamt__T_109_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_109_addr = 6'h27;
  assign queue_bits_wb_instr_shamt__T_109_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_109_en = reset;
  assign queue_bits_wb_instr_shamt__T_110_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_110_addr = 6'h28;
  assign queue_bits_wb_instr_shamt__T_110_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_110_en = reset;
  assign queue_bits_wb_instr_shamt__T_111_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_111_addr = 6'h29;
  assign queue_bits_wb_instr_shamt__T_111_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_111_en = reset;
  assign queue_bits_wb_instr_shamt__T_112_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_112_addr = 6'h2a;
  assign queue_bits_wb_instr_shamt__T_112_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_112_en = reset;
  assign queue_bits_wb_instr_shamt__T_113_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_113_addr = 6'h2b;
  assign queue_bits_wb_instr_shamt__T_113_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_113_en = reset;
  assign queue_bits_wb_instr_shamt__T_114_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_114_addr = 6'h2c;
  assign queue_bits_wb_instr_shamt__T_114_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_114_en = reset;
  assign queue_bits_wb_instr_shamt__T_115_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_115_addr = 6'h2d;
  assign queue_bits_wb_instr_shamt__T_115_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_115_en = reset;
  assign queue_bits_wb_instr_shamt__T_116_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_116_addr = 6'h2e;
  assign queue_bits_wb_instr_shamt__T_116_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_116_en = reset;
  assign queue_bits_wb_instr_shamt__T_117_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_117_addr = 6'h2f;
  assign queue_bits_wb_instr_shamt__T_117_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_117_en = reset;
  assign queue_bits_wb_instr_shamt__T_118_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_118_addr = 6'h30;
  assign queue_bits_wb_instr_shamt__T_118_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_118_en = reset;
  assign queue_bits_wb_instr_shamt__T_119_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_119_addr = 6'h31;
  assign queue_bits_wb_instr_shamt__T_119_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_119_en = reset;
  assign queue_bits_wb_instr_shamt__T_120_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_120_addr = 6'h32;
  assign queue_bits_wb_instr_shamt__T_120_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_120_en = reset;
  assign queue_bits_wb_instr_shamt__T_121_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_121_addr = 6'h33;
  assign queue_bits_wb_instr_shamt__T_121_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_121_en = reset;
  assign queue_bits_wb_instr_shamt__T_122_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_122_addr = 6'h34;
  assign queue_bits_wb_instr_shamt__T_122_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_122_en = reset;
  assign queue_bits_wb_instr_shamt__T_123_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_123_addr = 6'h35;
  assign queue_bits_wb_instr_shamt__T_123_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_123_en = reset;
  assign queue_bits_wb_instr_shamt__T_124_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_124_addr = 6'h36;
  assign queue_bits_wb_instr_shamt__T_124_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_124_en = reset;
  assign queue_bits_wb_instr_shamt__T_125_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_125_addr = 6'h37;
  assign queue_bits_wb_instr_shamt__T_125_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_125_en = reset;
  assign queue_bits_wb_instr_shamt__T_126_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_126_addr = 6'h38;
  assign queue_bits_wb_instr_shamt__T_126_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_126_en = reset;
  assign queue_bits_wb_instr_shamt__T_127_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_127_addr = 6'h39;
  assign queue_bits_wb_instr_shamt__T_127_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_127_en = reset;
  assign queue_bits_wb_instr_shamt__T_128_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_128_addr = 6'h3a;
  assign queue_bits_wb_instr_shamt__T_128_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_128_en = reset;
  assign queue_bits_wb_instr_shamt__T_129_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_129_addr = 6'h3b;
  assign queue_bits_wb_instr_shamt__T_129_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_129_en = reset;
  assign queue_bits_wb_instr_shamt__T_130_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_130_addr = 6'h3c;
  assign queue_bits_wb_instr_shamt__T_130_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_130_en = reset;
  assign queue_bits_wb_instr_shamt__T_131_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_131_addr = 6'h3d;
  assign queue_bits_wb_instr_shamt__T_131_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_131_en = reset;
  assign queue_bits_wb_instr_shamt__T_132_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_132_addr = 6'h3e;
  assign queue_bits_wb_instr_shamt__T_132_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_132_en = reset;
  assign queue_bits_wb_instr_shamt__T_133_data = 5'h0;
  assign queue_bits_wb_instr_shamt__T_133_addr = 6'h3f;
  assign queue_bits_wb_instr_shamt__T_133_mask = 1'h0;
  assign queue_bits_wb_instr_shamt__T_133_en = reset;
  assign queue_bits_wb_instr_shamt_q_head_w_data = 5'h0;
  assign queue_bits_wb_instr_shamt_q_head_w_addr = head;
  assign queue_bits_wb_instr_shamt_q_head_w_mask = 1'h0;
  assign queue_bits_wb_instr_shamt_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_instr_func_q_head_r_addr = head;
  assign queue_bits_wb_instr_func_q_head_r_data = queue_bits_wb_instr_func[queue_bits_wb_instr_func_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_instr_func__T_3_data = io_enq_0_bits_data_wb_instr_func;
  assign queue_bits_wb_instr_func__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_instr_func__T_3_mask = 1'h1;
  assign queue_bits_wb_instr_func__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_instr_func__T_4_data = io_enq_1_bits_data_wb_instr_func;
  assign queue_bits_wb_instr_func__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_instr_func__T_4_mask = 1'h1;
  assign queue_bits_wb_instr_func__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_instr_func__T_5_data = 6'h0;
  assign queue_bits_wb_instr_func__T_5_addr = 6'h0;
  assign queue_bits_wb_instr_func__T_5_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_5_en = 1'h0;
  assign queue_bits_wb_instr_func__T_6_data = 6'h0;
  assign queue_bits_wb_instr_func__T_6_addr = 6'h1;
  assign queue_bits_wb_instr_func__T_6_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_6_en = 1'h0;
  assign queue_bits_wb_instr_func__T_7_data = 6'h0;
  assign queue_bits_wb_instr_func__T_7_addr = 6'h2;
  assign queue_bits_wb_instr_func__T_7_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_7_en = 1'h0;
  assign queue_bits_wb_instr_func__T_8_data = 6'h0;
  assign queue_bits_wb_instr_func__T_8_addr = 6'h3;
  assign queue_bits_wb_instr_func__T_8_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_8_en = 1'h0;
  assign queue_bits_wb_instr_func__T_9_data = 6'h0;
  assign queue_bits_wb_instr_func__T_9_addr = 6'h4;
  assign queue_bits_wb_instr_func__T_9_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_9_en = 1'h0;
  assign queue_bits_wb_instr_func__T_10_data = 6'h0;
  assign queue_bits_wb_instr_func__T_10_addr = 6'h5;
  assign queue_bits_wb_instr_func__T_10_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_10_en = 1'h0;
  assign queue_bits_wb_instr_func__T_11_data = 6'h0;
  assign queue_bits_wb_instr_func__T_11_addr = 6'h6;
  assign queue_bits_wb_instr_func__T_11_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_11_en = 1'h0;
  assign queue_bits_wb_instr_func__T_12_data = 6'h0;
  assign queue_bits_wb_instr_func__T_12_addr = 6'h7;
  assign queue_bits_wb_instr_func__T_12_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_12_en = 1'h0;
  assign queue_bits_wb_instr_func__T_13_data = 6'h0;
  assign queue_bits_wb_instr_func__T_13_addr = 6'h8;
  assign queue_bits_wb_instr_func__T_13_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_13_en = 1'h0;
  assign queue_bits_wb_instr_func__T_14_data = 6'h0;
  assign queue_bits_wb_instr_func__T_14_addr = 6'h9;
  assign queue_bits_wb_instr_func__T_14_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_14_en = 1'h0;
  assign queue_bits_wb_instr_func__T_15_data = 6'h0;
  assign queue_bits_wb_instr_func__T_15_addr = 6'ha;
  assign queue_bits_wb_instr_func__T_15_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_15_en = 1'h0;
  assign queue_bits_wb_instr_func__T_16_data = 6'h0;
  assign queue_bits_wb_instr_func__T_16_addr = 6'hb;
  assign queue_bits_wb_instr_func__T_16_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_16_en = 1'h0;
  assign queue_bits_wb_instr_func__T_17_data = 6'h0;
  assign queue_bits_wb_instr_func__T_17_addr = 6'hc;
  assign queue_bits_wb_instr_func__T_17_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_17_en = 1'h0;
  assign queue_bits_wb_instr_func__T_18_data = 6'h0;
  assign queue_bits_wb_instr_func__T_18_addr = 6'hd;
  assign queue_bits_wb_instr_func__T_18_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_18_en = 1'h0;
  assign queue_bits_wb_instr_func__T_19_data = 6'h0;
  assign queue_bits_wb_instr_func__T_19_addr = 6'he;
  assign queue_bits_wb_instr_func__T_19_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_19_en = 1'h0;
  assign queue_bits_wb_instr_func__T_20_data = 6'h0;
  assign queue_bits_wb_instr_func__T_20_addr = 6'hf;
  assign queue_bits_wb_instr_func__T_20_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_20_en = 1'h0;
  assign queue_bits_wb_instr_func__T_21_data = 6'h0;
  assign queue_bits_wb_instr_func__T_21_addr = 6'h10;
  assign queue_bits_wb_instr_func__T_21_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_21_en = 1'h0;
  assign queue_bits_wb_instr_func__T_22_data = 6'h0;
  assign queue_bits_wb_instr_func__T_22_addr = 6'h11;
  assign queue_bits_wb_instr_func__T_22_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_22_en = 1'h0;
  assign queue_bits_wb_instr_func__T_23_data = 6'h0;
  assign queue_bits_wb_instr_func__T_23_addr = 6'h12;
  assign queue_bits_wb_instr_func__T_23_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_23_en = 1'h0;
  assign queue_bits_wb_instr_func__T_24_data = 6'h0;
  assign queue_bits_wb_instr_func__T_24_addr = 6'h13;
  assign queue_bits_wb_instr_func__T_24_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_24_en = 1'h0;
  assign queue_bits_wb_instr_func__T_25_data = 6'h0;
  assign queue_bits_wb_instr_func__T_25_addr = 6'h14;
  assign queue_bits_wb_instr_func__T_25_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_25_en = 1'h0;
  assign queue_bits_wb_instr_func__T_26_data = 6'h0;
  assign queue_bits_wb_instr_func__T_26_addr = 6'h15;
  assign queue_bits_wb_instr_func__T_26_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_26_en = 1'h0;
  assign queue_bits_wb_instr_func__T_27_data = 6'h0;
  assign queue_bits_wb_instr_func__T_27_addr = 6'h16;
  assign queue_bits_wb_instr_func__T_27_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_27_en = 1'h0;
  assign queue_bits_wb_instr_func__T_28_data = 6'h0;
  assign queue_bits_wb_instr_func__T_28_addr = 6'h17;
  assign queue_bits_wb_instr_func__T_28_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_28_en = 1'h0;
  assign queue_bits_wb_instr_func__T_29_data = 6'h0;
  assign queue_bits_wb_instr_func__T_29_addr = 6'h18;
  assign queue_bits_wb_instr_func__T_29_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_29_en = 1'h0;
  assign queue_bits_wb_instr_func__T_30_data = 6'h0;
  assign queue_bits_wb_instr_func__T_30_addr = 6'h19;
  assign queue_bits_wb_instr_func__T_30_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_30_en = 1'h0;
  assign queue_bits_wb_instr_func__T_31_data = 6'h0;
  assign queue_bits_wb_instr_func__T_31_addr = 6'h1a;
  assign queue_bits_wb_instr_func__T_31_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_31_en = 1'h0;
  assign queue_bits_wb_instr_func__T_32_data = 6'h0;
  assign queue_bits_wb_instr_func__T_32_addr = 6'h1b;
  assign queue_bits_wb_instr_func__T_32_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_32_en = 1'h0;
  assign queue_bits_wb_instr_func__T_33_data = 6'h0;
  assign queue_bits_wb_instr_func__T_33_addr = 6'h1c;
  assign queue_bits_wb_instr_func__T_33_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_33_en = 1'h0;
  assign queue_bits_wb_instr_func__T_34_data = 6'h0;
  assign queue_bits_wb_instr_func__T_34_addr = 6'h1d;
  assign queue_bits_wb_instr_func__T_34_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_34_en = 1'h0;
  assign queue_bits_wb_instr_func__T_35_data = 6'h0;
  assign queue_bits_wb_instr_func__T_35_addr = 6'h1e;
  assign queue_bits_wb_instr_func__T_35_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_35_en = 1'h0;
  assign queue_bits_wb_instr_func__T_36_data = 6'h0;
  assign queue_bits_wb_instr_func__T_36_addr = 6'h1f;
  assign queue_bits_wb_instr_func__T_36_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_36_en = 1'h0;
  assign queue_bits_wb_instr_func__T_37_data = 6'h0;
  assign queue_bits_wb_instr_func__T_37_addr = 6'h20;
  assign queue_bits_wb_instr_func__T_37_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_37_en = 1'h0;
  assign queue_bits_wb_instr_func__T_38_data = 6'h0;
  assign queue_bits_wb_instr_func__T_38_addr = 6'h21;
  assign queue_bits_wb_instr_func__T_38_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_38_en = 1'h0;
  assign queue_bits_wb_instr_func__T_39_data = 6'h0;
  assign queue_bits_wb_instr_func__T_39_addr = 6'h22;
  assign queue_bits_wb_instr_func__T_39_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_39_en = 1'h0;
  assign queue_bits_wb_instr_func__T_40_data = 6'h0;
  assign queue_bits_wb_instr_func__T_40_addr = 6'h23;
  assign queue_bits_wb_instr_func__T_40_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_40_en = 1'h0;
  assign queue_bits_wb_instr_func__T_41_data = 6'h0;
  assign queue_bits_wb_instr_func__T_41_addr = 6'h24;
  assign queue_bits_wb_instr_func__T_41_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_41_en = 1'h0;
  assign queue_bits_wb_instr_func__T_42_data = 6'h0;
  assign queue_bits_wb_instr_func__T_42_addr = 6'h25;
  assign queue_bits_wb_instr_func__T_42_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_42_en = 1'h0;
  assign queue_bits_wb_instr_func__T_43_data = 6'h0;
  assign queue_bits_wb_instr_func__T_43_addr = 6'h26;
  assign queue_bits_wb_instr_func__T_43_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_43_en = 1'h0;
  assign queue_bits_wb_instr_func__T_44_data = 6'h0;
  assign queue_bits_wb_instr_func__T_44_addr = 6'h27;
  assign queue_bits_wb_instr_func__T_44_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_44_en = 1'h0;
  assign queue_bits_wb_instr_func__T_45_data = 6'h0;
  assign queue_bits_wb_instr_func__T_45_addr = 6'h28;
  assign queue_bits_wb_instr_func__T_45_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_45_en = 1'h0;
  assign queue_bits_wb_instr_func__T_46_data = 6'h0;
  assign queue_bits_wb_instr_func__T_46_addr = 6'h29;
  assign queue_bits_wb_instr_func__T_46_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_46_en = 1'h0;
  assign queue_bits_wb_instr_func__T_47_data = 6'h0;
  assign queue_bits_wb_instr_func__T_47_addr = 6'h2a;
  assign queue_bits_wb_instr_func__T_47_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_47_en = 1'h0;
  assign queue_bits_wb_instr_func__T_48_data = 6'h0;
  assign queue_bits_wb_instr_func__T_48_addr = 6'h2b;
  assign queue_bits_wb_instr_func__T_48_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_48_en = 1'h0;
  assign queue_bits_wb_instr_func__T_49_data = 6'h0;
  assign queue_bits_wb_instr_func__T_49_addr = 6'h2c;
  assign queue_bits_wb_instr_func__T_49_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_49_en = 1'h0;
  assign queue_bits_wb_instr_func__T_50_data = 6'h0;
  assign queue_bits_wb_instr_func__T_50_addr = 6'h2d;
  assign queue_bits_wb_instr_func__T_50_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_50_en = 1'h0;
  assign queue_bits_wb_instr_func__T_51_data = 6'h0;
  assign queue_bits_wb_instr_func__T_51_addr = 6'h2e;
  assign queue_bits_wb_instr_func__T_51_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_51_en = 1'h0;
  assign queue_bits_wb_instr_func__T_52_data = 6'h0;
  assign queue_bits_wb_instr_func__T_52_addr = 6'h2f;
  assign queue_bits_wb_instr_func__T_52_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_52_en = 1'h0;
  assign queue_bits_wb_instr_func__T_53_data = 6'h0;
  assign queue_bits_wb_instr_func__T_53_addr = 6'h30;
  assign queue_bits_wb_instr_func__T_53_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_53_en = 1'h0;
  assign queue_bits_wb_instr_func__T_54_data = 6'h0;
  assign queue_bits_wb_instr_func__T_54_addr = 6'h31;
  assign queue_bits_wb_instr_func__T_54_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_54_en = 1'h0;
  assign queue_bits_wb_instr_func__T_55_data = 6'h0;
  assign queue_bits_wb_instr_func__T_55_addr = 6'h32;
  assign queue_bits_wb_instr_func__T_55_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_55_en = 1'h0;
  assign queue_bits_wb_instr_func__T_56_data = 6'h0;
  assign queue_bits_wb_instr_func__T_56_addr = 6'h33;
  assign queue_bits_wb_instr_func__T_56_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_56_en = 1'h0;
  assign queue_bits_wb_instr_func__T_57_data = 6'h0;
  assign queue_bits_wb_instr_func__T_57_addr = 6'h34;
  assign queue_bits_wb_instr_func__T_57_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_57_en = 1'h0;
  assign queue_bits_wb_instr_func__T_58_data = 6'h0;
  assign queue_bits_wb_instr_func__T_58_addr = 6'h35;
  assign queue_bits_wb_instr_func__T_58_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_58_en = 1'h0;
  assign queue_bits_wb_instr_func__T_59_data = 6'h0;
  assign queue_bits_wb_instr_func__T_59_addr = 6'h36;
  assign queue_bits_wb_instr_func__T_59_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_59_en = 1'h0;
  assign queue_bits_wb_instr_func__T_60_data = 6'h0;
  assign queue_bits_wb_instr_func__T_60_addr = 6'h37;
  assign queue_bits_wb_instr_func__T_60_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_60_en = 1'h0;
  assign queue_bits_wb_instr_func__T_61_data = 6'h0;
  assign queue_bits_wb_instr_func__T_61_addr = 6'h38;
  assign queue_bits_wb_instr_func__T_61_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_61_en = 1'h0;
  assign queue_bits_wb_instr_func__T_62_data = 6'h0;
  assign queue_bits_wb_instr_func__T_62_addr = 6'h39;
  assign queue_bits_wb_instr_func__T_62_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_62_en = 1'h0;
  assign queue_bits_wb_instr_func__T_63_data = 6'h0;
  assign queue_bits_wb_instr_func__T_63_addr = 6'h3a;
  assign queue_bits_wb_instr_func__T_63_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_63_en = 1'h0;
  assign queue_bits_wb_instr_func__T_64_data = 6'h0;
  assign queue_bits_wb_instr_func__T_64_addr = 6'h3b;
  assign queue_bits_wb_instr_func__T_64_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_64_en = 1'h0;
  assign queue_bits_wb_instr_func__T_65_data = 6'h0;
  assign queue_bits_wb_instr_func__T_65_addr = 6'h3c;
  assign queue_bits_wb_instr_func__T_65_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_65_en = 1'h0;
  assign queue_bits_wb_instr_func__T_66_data = 6'h0;
  assign queue_bits_wb_instr_func__T_66_addr = 6'h3d;
  assign queue_bits_wb_instr_func__T_66_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_66_en = 1'h0;
  assign queue_bits_wb_instr_func__T_67_data = 6'h0;
  assign queue_bits_wb_instr_func__T_67_addr = 6'h3e;
  assign queue_bits_wb_instr_func__T_67_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_67_en = 1'h0;
  assign queue_bits_wb_instr_func__T_68_data = 6'h0;
  assign queue_bits_wb_instr_func__T_68_addr = 6'h3f;
  assign queue_bits_wb_instr_func__T_68_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_68_en = 1'h0;
  assign queue_bits_wb_instr_func__T_70_data = 6'h0;
  assign queue_bits_wb_instr_func__T_70_addr = 6'h0;
  assign queue_bits_wb_instr_func__T_70_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_70_en = reset;
  assign queue_bits_wb_instr_func__T_71_data = 6'h0;
  assign queue_bits_wb_instr_func__T_71_addr = 6'h1;
  assign queue_bits_wb_instr_func__T_71_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_71_en = reset;
  assign queue_bits_wb_instr_func__T_72_data = 6'h0;
  assign queue_bits_wb_instr_func__T_72_addr = 6'h2;
  assign queue_bits_wb_instr_func__T_72_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_72_en = reset;
  assign queue_bits_wb_instr_func__T_73_data = 6'h0;
  assign queue_bits_wb_instr_func__T_73_addr = 6'h3;
  assign queue_bits_wb_instr_func__T_73_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_73_en = reset;
  assign queue_bits_wb_instr_func__T_74_data = 6'h0;
  assign queue_bits_wb_instr_func__T_74_addr = 6'h4;
  assign queue_bits_wb_instr_func__T_74_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_74_en = reset;
  assign queue_bits_wb_instr_func__T_75_data = 6'h0;
  assign queue_bits_wb_instr_func__T_75_addr = 6'h5;
  assign queue_bits_wb_instr_func__T_75_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_75_en = reset;
  assign queue_bits_wb_instr_func__T_76_data = 6'h0;
  assign queue_bits_wb_instr_func__T_76_addr = 6'h6;
  assign queue_bits_wb_instr_func__T_76_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_76_en = reset;
  assign queue_bits_wb_instr_func__T_77_data = 6'h0;
  assign queue_bits_wb_instr_func__T_77_addr = 6'h7;
  assign queue_bits_wb_instr_func__T_77_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_77_en = reset;
  assign queue_bits_wb_instr_func__T_78_data = 6'h0;
  assign queue_bits_wb_instr_func__T_78_addr = 6'h8;
  assign queue_bits_wb_instr_func__T_78_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_78_en = reset;
  assign queue_bits_wb_instr_func__T_79_data = 6'h0;
  assign queue_bits_wb_instr_func__T_79_addr = 6'h9;
  assign queue_bits_wb_instr_func__T_79_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_79_en = reset;
  assign queue_bits_wb_instr_func__T_80_data = 6'h0;
  assign queue_bits_wb_instr_func__T_80_addr = 6'ha;
  assign queue_bits_wb_instr_func__T_80_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_80_en = reset;
  assign queue_bits_wb_instr_func__T_81_data = 6'h0;
  assign queue_bits_wb_instr_func__T_81_addr = 6'hb;
  assign queue_bits_wb_instr_func__T_81_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_81_en = reset;
  assign queue_bits_wb_instr_func__T_82_data = 6'h0;
  assign queue_bits_wb_instr_func__T_82_addr = 6'hc;
  assign queue_bits_wb_instr_func__T_82_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_82_en = reset;
  assign queue_bits_wb_instr_func__T_83_data = 6'h0;
  assign queue_bits_wb_instr_func__T_83_addr = 6'hd;
  assign queue_bits_wb_instr_func__T_83_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_83_en = reset;
  assign queue_bits_wb_instr_func__T_84_data = 6'h0;
  assign queue_bits_wb_instr_func__T_84_addr = 6'he;
  assign queue_bits_wb_instr_func__T_84_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_84_en = reset;
  assign queue_bits_wb_instr_func__T_85_data = 6'h0;
  assign queue_bits_wb_instr_func__T_85_addr = 6'hf;
  assign queue_bits_wb_instr_func__T_85_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_85_en = reset;
  assign queue_bits_wb_instr_func__T_86_data = 6'h0;
  assign queue_bits_wb_instr_func__T_86_addr = 6'h10;
  assign queue_bits_wb_instr_func__T_86_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_86_en = reset;
  assign queue_bits_wb_instr_func__T_87_data = 6'h0;
  assign queue_bits_wb_instr_func__T_87_addr = 6'h11;
  assign queue_bits_wb_instr_func__T_87_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_87_en = reset;
  assign queue_bits_wb_instr_func__T_88_data = 6'h0;
  assign queue_bits_wb_instr_func__T_88_addr = 6'h12;
  assign queue_bits_wb_instr_func__T_88_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_88_en = reset;
  assign queue_bits_wb_instr_func__T_89_data = 6'h0;
  assign queue_bits_wb_instr_func__T_89_addr = 6'h13;
  assign queue_bits_wb_instr_func__T_89_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_89_en = reset;
  assign queue_bits_wb_instr_func__T_90_data = 6'h0;
  assign queue_bits_wb_instr_func__T_90_addr = 6'h14;
  assign queue_bits_wb_instr_func__T_90_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_90_en = reset;
  assign queue_bits_wb_instr_func__T_91_data = 6'h0;
  assign queue_bits_wb_instr_func__T_91_addr = 6'h15;
  assign queue_bits_wb_instr_func__T_91_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_91_en = reset;
  assign queue_bits_wb_instr_func__T_92_data = 6'h0;
  assign queue_bits_wb_instr_func__T_92_addr = 6'h16;
  assign queue_bits_wb_instr_func__T_92_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_92_en = reset;
  assign queue_bits_wb_instr_func__T_93_data = 6'h0;
  assign queue_bits_wb_instr_func__T_93_addr = 6'h17;
  assign queue_bits_wb_instr_func__T_93_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_93_en = reset;
  assign queue_bits_wb_instr_func__T_94_data = 6'h0;
  assign queue_bits_wb_instr_func__T_94_addr = 6'h18;
  assign queue_bits_wb_instr_func__T_94_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_94_en = reset;
  assign queue_bits_wb_instr_func__T_95_data = 6'h0;
  assign queue_bits_wb_instr_func__T_95_addr = 6'h19;
  assign queue_bits_wb_instr_func__T_95_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_95_en = reset;
  assign queue_bits_wb_instr_func__T_96_data = 6'h0;
  assign queue_bits_wb_instr_func__T_96_addr = 6'h1a;
  assign queue_bits_wb_instr_func__T_96_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_96_en = reset;
  assign queue_bits_wb_instr_func__T_97_data = 6'h0;
  assign queue_bits_wb_instr_func__T_97_addr = 6'h1b;
  assign queue_bits_wb_instr_func__T_97_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_97_en = reset;
  assign queue_bits_wb_instr_func__T_98_data = 6'h0;
  assign queue_bits_wb_instr_func__T_98_addr = 6'h1c;
  assign queue_bits_wb_instr_func__T_98_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_98_en = reset;
  assign queue_bits_wb_instr_func__T_99_data = 6'h0;
  assign queue_bits_wb_instr_func__T_99_addr = 6'h1d;
  assign queue_bits_wb_instr_func__T_99_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_99_en = reset;
  assign queue_bits_wb_instr_func__T_100_data = 6'h0;
  assign queue_bits_wb_instr_func__T_100_addr = 6'h1e;
  assign queue_bits_wb_instr_func__T_100_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_100_en = reset;
  assign queue_bits_wb_instr_func__T_101_data = 6'h0;
  assign queue_bits_wb_instr_func__T_101_addr = 6'h1f;
  assign queue_bits_wb_instr_func__T_101_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_101_en = reset;
  assign queue_bits_wb_instr_func__T_102_data = 6'h0;
  assign queue_bits_wb_instr_func__T_102_addr = 6'h20;
  assign queue_bits_wb_instr_func__T_102_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_102_en = reset;
  assign queue_bits_wb_instr_func__T_103_data = 6'h0;
  assign queue_bits_wb_instr_func__T_103_addr = 6'h21;
  assign queue_bits_wb_instr_func__T_103_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_103_en = reset;
  assign queue_bits_wb_instr_func__T_104_data = 6'h0;
  assign queue_bits_wb_instr_func__T_104_addr = 6'h22;
  assign queue_bits_wb_instr_func__T_104_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_104_en = reset;
  assign queue_bits_wb_instr_func__T_105_data = 6'h0;
  assign queue_bits_wb_instr_func__T_105_addr = 6'h23;
  assign queue_bits_wb_instr_func__T_105_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_105_en = reset;
  assign queue_bits_wb_instr_func__T_106_data = 6'h0;
  assign queue_bits_wb_instr_func__T_106_addr = 6'h24;
  assign queue_bits_wb_instr_func__T_106_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_106_en = reset;
  assign queue_bits_wb_instr_func__T_107_data = 6'h0;
  assign queue_bits_wb_instr_func__T_107_addr = 6'h25;
  assign queue_bits_wb_instr_func__T_107_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_107_en = reset;
  assign queue_bits_wb_instr_func__T_108_data = 6'h0;
  assign queue_bits_wb_instr_func__T_108_addr = 6'h26;
  assign queue_bits_wb_instr_func__T_108_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_108_en = reset;
  assign queue_bits_wb_instr_func__T_109_data = 6'h0;
  assign queue_bits_wb_instr_func__T_109_addr = 6'h27;
  assign queue_bits_wb_instr_func__T_109_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_109_en = reset;
  assign queue_bits_wb_instr_func__T_110_data = 6'h0;
  assign queue_bits_wb_instr_func__T_110_addr = 6'h28;
  assign queue_bits_wb_instr_func__T_110_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_110_en = reset;
  assign queue_bits_wb_instr_func__T_111_data = 6'h0;
  assign queue_bits_wb_instr_func__T_111_addr = 6'h29;
  assign queue_bits_wb_instr_func__T_111_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_111_en = reset;
  assign queue_bits_wb_instr_func__T_112_data = 6'h0;
  assign queue_bits_wb_instr_func__T_112_addr = 6'h2a;
  assign queue_bits_wb_instr_func__T_112_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_112_en = reset;
  assign queue_bits_wb_instr_func__T_113_data = 6'h0;
  assign queue_bits_wb_instr_func__T_113_addr = 6'h2b;
  assign queue_bits_wb_instr_func__T_113_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_113_en = reset;
  assign queue_bits_wb_instr_func__T_114_data = 6'h0;
  assign queue_bits_wb_instr_func__T_114_addr = 6'h2c;
  assign queue_bits_wb_instr_func__T_114_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_114_en = reset;
  assign queue_bits_wb_instr_func__T_115_data = 6'h0;
  assign queue_bits_wb_instr_func__T_115_addr = 6'h2d;
  assign queue_bits_wb_instr_func__T_115_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_115_en = reset;
  assign queue_bits_wb_instr_func__T_116_data = 6'h0;
  assign queue_bits_wb_instr_func__T_116_addr = 6'h2e;
  assign queue_bits_wb_instr_func__T_116_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_116_en = reset;
  assign queue_bits_wb_instr_func__T_117_data = 6'h0;
  assign queue_bits_wb_instr_func__T_117_addr = 6'h2f;
  assign queue_bits_wb_instr_func__T_117_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_117_en = reset;
  assign queue_bits_wb_instr_func__T_118_data = 6'h0;
  assign queue_bits_wb_instr_func__T_118_addr = 6'h30;
  assign queue_bits_wb_instr_func__T_118_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_118_en = reset;
  assign queue_bits_wb_instr_func__T_119_data = 6'h0;
  assign queue_bits_wb_instr_func__T_119_addr = 6'h31;
  assign queue_bits_wb_instr_func__T_119_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_119_en = reset;
  assign queue_bits_wb_instr_func__T_120_data = 6'h0;
  assign queue_bits_wb_instr_func__T_120_addr = 6'h32;
  assign queue_bits_wb_instr_func__T_120_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_120_en = reset;
  assign queue_bits_wb_instr_func__T_121_data = 6'h0;
  assign queue_bits_wb_instr_func__T_121_addr = 6'h33;
  assign queue_bits_wb_instr_func__T_121_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_121_en = reset;
  assign queue_bits_wb_instr_func__T_122_data = 6'h0;
  assign queue_bits_wb_instr_func__T_122_addr = 6'h34;
  assign queue_bits_wb_instr_func__T_122_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_122_en = reset;
  assign queue_bits_wb_instr_func__T_123_data = 6'h0;
  assign queue_bits_wb_instr_func__T_123_addr = 6'h35;
  assign queue_bits_wb_instr_func__T_123_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_123_en = reset;
  assign queue_bits_wb_instr_func__T_124_data = 6'h0;
  assign queue_bits_wb_instr_func__T_124_addr = 6'h36;
  assign queue_bits_wb_instr_func__T_124_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_124_en = reset;
  assign queue_bits_wb_instr_func__T_125_data = 6'h0;
  assign queue_bits_wb_instr_func__T_125_addr = 6'h37;
  assign queue_bits_wb_instr_func__T_125_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_125_en = reset;
  assign queue_bits_wb_instr_func__T_126_data = 6'h0;
  assign queue_bits_wb_instr_func__T_126_addr = 6'h38;
  assign queue_bits_wb_instr_func__T_126_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_126_en = reset;
  assign queue_bits_wb_instr_func__T_127_data = 6'h0;
  assign queue_bits_wb_instr_func__T_127_addr = 6'h39;
  assign queue_bits_wb_instr_func__T_127_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_127_en = reset;
  assign queue_bits_wb_instr_func__T_128_data = 6'h0;
  assign queue_bits_wb_instr_func__T_128_addr = 6'h3a;
  assign queue_bits_wb_instr_func__T_128_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_128_en = reset;
  assign queue_bits_wb_instr_func__T_129_data = 6'h0;
  assign queue_bits_wb_instr_func__T_129_addr = 6'h3b;
  assign queue_bits_wb_instr_func__T_129_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_129_en = reset;
  assign queue_bits_wb_instr_func__T_130_data = 6'h0;
  assign queue_bits_wb_instr_func__T_130_addr = 6'h3c;
  assign queue_bits_wb_instr_func__T_130_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_130_en = reset;
  assign queue_bits_wb_instr_func__T_131_data = 6'h0;
  assign queue_bits_wb_instr_func__T_131_addr = 6'h3d;
  assign queue_bits_wb_instr_func__T_131_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_131_en = reset;
  assign queue_bits_wb_instr_func__T_132_data = 6'h0;
  assign queue_bits_wb_instr_func__T_132_addr = 6'h3e;
  assign queue_bits_wb_instr_func__T_132_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_132_en = reset;
  assign queue_bits_wb_instr_func__T_133_data = 6'h0;
  assign queue_bits_wb_instr_func__T_133_addr = 6'h3f;
  assign queue_bits_wb_instr_func__T_133_mask = 1'h0;
  assign queue_bits_wb_instr_func__T_133_en = reset;
  assign queue_bits_wb_instr_func_q_head_w_data = 6'h0;
  assign queue_bits_wb_instr_func_q_head_w_addr = head;
  assign queue_bits_wb_instr_func_q_head_w_mask = 1'h0;
  assign queue_bits_wb_instr_func_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_rd_idx_q_head_r_addr = head;
  assign queue_bits_wb_rd_idx_q_head_r_data = queue_bits_wb_rd_idx[queue_bits_wb_rd_idx_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_rd_idx__T_3_data = io_enq_0_bits_data_wb_rd_idx;
  assign queue_bits_wb_rd_idx__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_rd_idx__T_3_mask = 1'h1;
  assign queue_bits_wb_rd_idx__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_rd_idx__T_4_data = io_enq_1_bits_data_wb_rd_idx;
  assign queue_bits_wb_rd_idx__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_rd_idx__T_4_mask = 1'h1;
  assign queue_bits_wb_rd_idx__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_rd_idx__T_5_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_5_addr = 6'h0;
  assign queue_bits_wb_rd_idx__T_5_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_5_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_6_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_6_addr = 6'h1;
  assign queue_bits_wb_rd_idx__T_6_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_6_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_7_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_7_addr = 6'h2;
  assign queue_bits_wb_rd_idx__T_7_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_7_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_8_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_8_addr = 6'h3;
  assign queue_bits_wb_rd_idx__T_8_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_8_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_9_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_9_addr = 6'h4;
  assign queue_bits_wb_rd_idx__T_9_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_9_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_10_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_10_addr = 6'h5;
  assign queue_bits_wb_rd_idx__T_10_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_10_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_11_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_11_addr = 6'h6;
  assign queue_bits_wb_rd_idx__T_11_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_11_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_12_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_12_addr = 6'h7;
  assign queue_bits_wb_rd_idx__T_12_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_12_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_13_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_13_addr = 6'h8;
  assign queue_bits_wb_rd_idx__T_13_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_13_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_14_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_14_addr = 6'h9;
  assign queue_bits_wb_rd_idx__T_14_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_14_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_15_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_15_addr = 6'ha;
  assign queue_bits_wb_rd_idx__T_15_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_15_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_16_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_16_addr = 6'hb;
  assign queue_bits_wb_rd_idx__T_16_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_16_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_17_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_17_addr = 6'hc;
  assign queue_bits_wb_rd_idx__T_17_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_17_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_18_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_18_addr = 6'hd;
  assign queue_bits_wb_rd_idx__T_18_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_18_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_19_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_19_addr = 6'he;
  assign queue_bits_wb_rd_idx__T_19_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_19_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_20_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_20_addr = 6'hf;
  assign queue_bits_wb_rd_idx__T_20_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_20_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_21_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_21_addr = 6'h10;
  assign queue_bits_wb_rd_idx__T_21_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_21_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_22_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_22_addr = 6'h11;
  assign queue_bits_wb_rd_idx__T_22_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_22_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_23_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_23_addr = 6'h12;
  assign queue_bits_wb_rd_idx__T_23_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_23_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_24_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_24_addr = 6'h13;
  assign queue_bits_wb_rd_idx__T_24_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_24_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_25_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_25_addr = 6'h14;
  assign queue_bits_wb_rd_idx__T_25_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_25_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_26_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_26_addr = 6'h15;
  assign queue_bits_wb_rd_idx__T_26_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_26_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_27_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_27_addr = 6'h16;
  assign queue_bits_wb_rd_idx__T_27_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_27_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_28_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_28_addr = 6'h17;
  assign queue_bits_wb_rd_idx__T_28_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_28_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_29_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_29_addr = 6'h18;
  assign queue_bits_wb_rd_idx__T_29_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_29_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_30_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_30_addr = 6'h19;
  assign queue_bits_wb_rd_idx__T_30_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_30_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_31_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_31_addr = 6'h1a;
  assign queue_bits_wb_rd_idx__T_31_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_31_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_32_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_32_addr = 6'h1b;
  assign queue_bits_wb_rd_idx__T_32_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_32_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_33_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_33_addr = 6'h1c;
  assign queue_bits_wb_rd_idx__T_33_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_33_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_34_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_34_addr = 6'h1d;
  assign queue_bits_wb_rd_idx__T_34_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_34_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_35_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_35_addr = 6'h1e;
  assign queue_bits_wb_rd_idx__T_35_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_35_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_36_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_36_addr = 6'h1f;
  assign queue_bits_wb_rd_idx__T_36_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_36_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_37_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_37_addr = 6'h20;
  assign queue_bits_wb_rd_idx__T_37_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_37_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_38_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_38_addr = 6'h21;
  assign queue_bits_wb_rd_idx__T_38_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_38_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_39_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_39_addr = 6'h22;
  assign queue_bits_wb_rd_idx__T_39_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_39_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_40_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_40_addr = 6'h23;
  assign queue_bits_wb_rd_idx__T_40_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_40_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_41_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_41_addr = 6'h24;
  assign queue_bits_wb_rd_idx__T_41_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_41_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_42_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_42_addr = 6'h25;
  assign queue_bits_wb_rd_idx__T_42_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_42_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_43_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_43_addr = 6'h26;
  assign queue_bits_wb_rd_idx__T_43_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_43_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_44_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_44_addr = 6'h27;
  assign queue_bits_wb_rd_idx__T_44_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_44_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_45_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_45_addr = 6'h28;
  assign queue_bits_wb_rd_idx__T_45_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_45_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_46_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_46_addr = 6'h29;
  assign queue_bits_wb_rd_idx__T_46_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_46_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_47_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_47_addr = 6'h2a;
  assign queue_bits_wb_rd_idx__T_47_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_47_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_48_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_48_addr = 6'h2b;
  assign queue_bits_wb_rd_idx__T_48_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_48_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_49_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_49_addr = 6'h2c;
  assign queue_bits_wb_rd_idx__T_49_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_49_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_50_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_50_addr = 6'h2d;
  assign queue_bits_wb_rd_idx__T_50_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_50_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_51_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_51_addr = 6'h2e;
  assign queue_bits_wb_rd_idx__T_51_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_51_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_52_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_52_addr = 6'h2f;
  assign queue_bits_wb_rd_idx__T_52_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_52_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_53_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_53_addr = 6'h30;
  assign queue_bits_wb_rd_idx__T_53_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_53_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_54_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_54_addr = 6'h31;
  assign queue_bits_wb_rd_idx__T_54_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_54_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_55_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_55_addr = 6'h32;
  assign queue_bits_wb_rd_idx__T_55_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_55_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_56_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_56_addr = 6'h33;
  assign queue_bits_wb_rd_idx__T_56_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_56_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_57_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_57_addr = 6'h34;
  assign queue_bits_wb_rd_idx__T_57_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_57_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_58_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_58_addr = 6'h35;
  assign queue_bits_wb_rd_idx__T_58_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_58_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_59_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_59_addr = 6'h36;
  assign queue_bits_wb_rd_idx__T_59_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_59_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_60_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_60_addr = 6'h37;
  assign queue_bits_wb_rd_idx__T_60_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_60_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_61_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_61_addr = 6'h38;
  assign queue_bits_wb_rd_idx__T_61_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_61_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_62_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_62_addr = 6'h39;
  assign queue_bits_wb_rd_idx__T_62_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_62_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_63_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_63_addr = 6'h3a;
  assign queue_bits_wb_rd_idx__T_63_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_63_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_64_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_64_addr = 6'h3b;
  assign queue_bits_wb_rd_idx__T_64_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_64_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_65_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_65_addr = 6'h3c;
  assign queue_bits_wb_rd_idx__T_65_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_65_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_66_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_66_addr = 6'h3d;
  assign queue_bits_wb_rd_idx__T_66_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_66_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_67_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_67_addr = 6'h3e;
  assign queue_bits_wb_rd_idx__T_67_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_67_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_68_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_68_addr = 6'h3f;
  assign queue_bits_wb_rd_idx__T_68_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_68_en = 1'h0;
  assign queue_bits_wb_rd_idx__T_70_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_70_addr = 6'h0;
  assign queue_bits_wb_rd_idx__T_70_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_70_en = reset;
  assign queue_bits_wb_rd_idx__T_71_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_71_addr = 6'h1;
  assign queue_bits_wb_rd_idx__T_71_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_71_en = reset;
  assign queue_bits_wb_rd_idx__T_72_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_72_addr = 6'h2;
  assign queue_bits_wb_rd_idx__T_72_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_72_en = reset;
  assign queue_bits_wb_rd_idx__T_73_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_73_addr = 6'h3;
  assign queue_bits_wb_rd_idx__T_73_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_73_en = reset;
  assign queue_bits_wb_rd_idx__T_74_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_74_addr = 6'h4;
  assign queue_bits_wb_rd_idx__T_74_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_74_en = reset;
  assign queue_bits_wb_rd_idx__T_75_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_75_addr = 6'h5;
  assign queue_bits_wb_rd_idx__T_75_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_75_en = reset;
  assign queue_bits_wb_rd_idx__T_76_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_76_addr = 6'h6;
  assign queue_bits_wb_rd_idx__T_76_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_76_en = reset;
  assign queue_bits_wb_rd_idx__T_77_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_77_addr = 6'h7;
  assign queue_bits_wb_rd_idx__T_77_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_77_en = reset;
  assign queue_bits_wb_rd_idx__T_78_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_78_addr = 6'h8;
  assign queue_bits_wb_rd_idx__T_78_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_78_en = reset;
  assign queue_bits_wb_rd_idx__T_79_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_79_addr = 6'h9;
  assign queue_bits_wb_rd_idx__T_79_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_79_en = reset;
  assign queue_bits_wb_rd_idx__T_80_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_80_addr = 6'ha;
  assign queue_bits_wb_rd_idx__T_80_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_80_en = reset;
  assign queue_bits_wb_rd_idx__T_81_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_81_addr = 6'hb;
  assign queue_bits_wb_rd_idx__T_81_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_81_en = reset;
  assign queue_bits_wb_rd_idx__T_82_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_82_addr = 6'hc;
  assign queue_bits_wb_rd_idx__T_82_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_82_en = reset;
  assign queue_bits_wb_rd_idx__T_83_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_83_addr = 6'hd;
  assign queue_bits_wb_rd_idx__T_83_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_83_en = reset;
  assign queue_bits_wb_rd_idx__T_84_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_84_addr = 6'he;
  assign queue_bits_wb_rd_idx__T_84_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_84_en = reset;
  assign queue_bits_wb_rd_idx__T_85_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_85_addr = 6'hf;
  assign queue_bits_wb_rd_idx__T_85_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_85_en = reset;
  assign queue_bits_wb_rd_idx__T_86_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_86_addr = 6'h10;
  assign queue_bits_wb_rd_idx__T_86_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_86_en = reset;
  assign queue_bits_wb_rd_idx__T_87_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_87_addr = 6'h11;
  assign queue_bits_wb_rd_idx__T_87_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_87_en = reset;
  assign queue_bits_wb_rd_idx__T_88_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_88_addr = 6'h12;
  assign queue_bits_wb_rd_idx__T_88_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_88_en = reset;
  assign queue_bits_wb_rd_idx__T_89_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_89_addr = 6'h13;
  assign queue_bits_wb_rd_idx__T_89_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_89_en = reset;
  assign queue_bits_wb_rd_idx__T_90_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_90_addr = 6'h14;
  assign queue_bits_wb_rd_idx__T_90_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_90_en = reset;
  assign queue_bits_wb_rd_idx__T_91_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_91_addr = 6'h15;
  assign queue_bits_wb_rd_idx__T_91_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_91_en = reset;
  assign queue_bits_wb_rd_idx__T_92_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_92_addr = 6'h16;
  assign queue_bits_wb_rd_idx__T_92_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_92_en = reset;
  assign queue_bits_wb_rd_idx__T_93_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_93_addr = 6'h17;
  assign queue_bits_wb_rd_idx__T_93_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_93_en = reset;
  assign queue_bits_wb_rd_idx__T_94_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_94_addr = 6'h18;
  assign queue_bits_wb_rd_idx__T_94_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_94_en = reset;
  assign queue_bits_wb_rd_idx__T_95_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_95_addr = 6'h19;
  assign queue_bits_wb_rd_idx__T_95_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_95_en = reset;
  assign queue_bits_wb_rd_idx__T_96_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_96_addr = 6'h1a;
  assign queue_bits_wb_rd_idx__T_96_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_96_en = reset;
  assign queue_bits_wb_rd_idx__T_97_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_97_addr = 6'h1b;
  assign queue_bits_wb_rd_idx__T_97_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_97_en = reset;
  assign queue_bits_wb_rd_idx__T_98_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_98_addr = 6'h1c;
  assign queue_bits_wb_rd_idx__T_98_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_98_en = reset;
  assign queue_bits_wb_rd_idx__T_99_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_99_addr = 6'h1d;
  assign queue_bits_wb_rd_idx__T_99_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_99_en = reset;
  assign queue_bits_wb_rd_idx__T_100_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_100_addr = 6'h1e;
  assign queue_bits_wb_rd_idx__T_100_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_100_en = reset;
  assign queue_bits_wb_rd_idx__T_101_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_101_addr = 6'h1f;
  assign queue_bits_wb_rd_idx__T_101_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_101_en = reset;
  assign queue_bits_wb_rd_idx__T_102_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_102_addr = 6'h20;
  assign queue_bits_wb_rd_idx__T_102_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_102_en = reset;
  assign queue_bits_wb_rd_idx__T_103_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_103_addr = 6'h21;
  assign queue_bits_wb_rd_idx__T_103_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_103_en = reset;
  assign queue_bits_wb_rd_idx__T_104_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_104_addr = 6'h22;
  assign queue_bits_wb_rd_idx__T_104_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_104_en = reset;
  assign queue_bits_wb_rd_idx__T_105_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_105_addr = 6'h23;
  assign queue_bits_wb_rd_idx__T_105_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_105_en = reset;
  assign queue_bits_wb_rd_idx__T_106_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_106_addr = 6'h24;
  assign queue_bits_wb_rd_idx__T_106_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_106_en = reset;
  assign queue_bits_wb_rd_idx__T_107_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_107_addr = 6'h25;
  assign queue_bits_wb_rd_idx__T_107_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_107_en = reset;
  assign queue_bits_wb_rd_idx__T_108_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_108_addr = 6'h26;
  assign queue_bits_wb_rd_idx__T_108_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_108_en = reset;
  assign queue_bits_wb_rd_idx__T_109_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_109_addr = 6'h27;
  assign queue_bits_wb_rd_idx__T_109_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_109_en = reset;
  assign queue_bits_wb_rd_idx__T_110_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_110_addr = 6'h28;
  assign queue_bits_wb_rd_idx__T_110_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_110_en = reset;
  assign queue_bits_wb_rd_idx__T_111_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_111_addr = 6'h29;
  assign queue_bits_wb_rd_idx__T_111_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_111_en = reset;
  assign queue_bits_wb_rd_idx__T_112_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_112_addr = 6'h2a;
  assign queue_bits_wb_rd_idx__T_112_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_112_en = reset;
  assign queue_bits_wb_rd_idx__T_113_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_113_addr = 6'h2b;
  assign queue_bits_wb_rd_idx__T_113_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_113_en = reset;
  assign queue_bits_wb_rd_idx__T_114_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_114_addr = 6'h2c;
  assign queue_bits_wb_rd_idx__T_114_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_114_en = reset;
  assign queue_bits_wb_rd_idx__T_115_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_115_addr = 6'h2d;
  assign queue_bits_wb_rd_idx__T_115_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_115_en = reset;
  assign queue_bits_wb_rd_idx__T_116_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_116_addr = 6'h2e;
  assign queue_bits_wb_rd_idx__T_116_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_116_en = reset;
  assign queue_bits_wb_rd_idx__T_117_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_117_addr = 6'h2f;
  assign queue_bits_wb_rd_idx__T_117_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_117_en = reset;
  assign queue_bits_wb_rd_idx__T_118_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_118_addr = 6'h30;
  assign queue_bits_wb_rd_idx__T_118_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_118_en = reset;
  assign queue_bits_wb_rd_idx__T_119_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_119_addr = 6'h31;
  assign queue_bits_wb_rd_idx__T_119_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_119_en = reset;
  assign queue_bits_wb_rd_idx__T_120_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_120_addr = 6'h32;
  assign queue_bits_wb_rd_idx__T_120_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_120_en = reset;
  assign queue_bits_wb_rd_idx__T_121_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_121_addr = 6'h33;
  assign queue_bits_wb_rd_idx__T_121_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_121_en = reset;
  assign queue_bits_wb_rd_idx__T_122_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_122_addr = 6'h34;
  assign queue_bits_wb_rd_idx__T_122_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_122_en = reset;
  assign queue_bits_wb_rd_idx__T_123_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_123_addr = 6'h35;
  assign queue_bits_wb_rd_idx__T_123_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_123_en = reset;
  assign queue_bits_wb_rd_idx__T_124_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_124_addr = 6'h36;
  assign queue_bits_wb_rd_idx__T_124_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_124_en = reset;
  assign queue_bits_wb_rd_idx__T_125_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_125_addr = 6'h37;
  assign queue_bits_wb_rd_idx__T_125_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_125_en = reset;
  assign queue_bits_wb_rd_idx__T_126_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_126_addr = 6'h38;
  assign queue_bits_wb_rd_idx__T_126_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_126_en = reset;
  assign queue_bits_wb_rd_idx__T_127_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_127_addr = 6'h39;
  assign queue_bits_wb_rd_idx__T_127_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_127_en = reset;
  assign queue_bits_wb_rd_idx__T_128_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_128_addr = 6'h3a;
  assign queue_bits_wb_rd_idx__T_128_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_128_en = reset;
  assign queue_bits_wb_rd_idx__T_129_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_129_addr = 6'h3b;
  assign queue_bits_wb_rd_idx__T_129_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_129_en = reset;
  assign queue_bits_wb_rd_idx__T_130_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_130_addr = 6'h3c;
  assign queue_bits_wb_rd_idx__T_130_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_130_en = reset;
  assign queue_bits_wb_rd_idx__T_131_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_131_addr = 6'h3d;
  assign queue_bits_wb_rd_idx__T_131_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_131_en = reset;
  assign queue_bits_wb_rd_idx__T_132_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_132_addr = 6'h3e;
  assign queue_bits_wb_rd_idx__T_132_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_132_en = reset;
  assign queue_bits_wb_rd_idx__T_133_data = 5'h0;
  assign queue_bits_wb_rd_idx__T_133_addr = 6'h3f;
  assign queue_bits_wb_rd_idx__T_133_mask = 1'h0;
  assign queue_bits_wb_rd_idx__T_133_en = reset;
  assign queue_bits_wb_rd_idx_q_head_w_data = 5'h0;
  assign queue_bits_wb_rd_idx_q_head_w_addr = head;
  assign queue_bits_wb_rd_idx_q_head_w_mask = 1'h0;
  assign queue_bits_wb_rd_idx_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_ip7_q_head_r_addr = head;
  assign queue_bits_wb_ip7_q_head_r_data = queue_bits_wb_ip7[queue_bits_wb_ip7_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_ip7__T_3_data = io_enq_0_bits_data_wb_ip7;
  assign queue_bits_wb_ip7__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_ip7__T_3_mask = 1'h1;
  assign queue_bits_wb_ip7__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_ip7__T_4_data = io_enq_1_bits_data_wb_ip7;
  assign queue_bits_wb_ip7__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_ip7__T_4_mask = 1'h1;
  assign queue_bits_wb_ip7__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_ip7__T_5_data = 1'h0;
  assign queue_bits_wb_ip7__T_5_addr = 6'h0;
  assign queue_bits_wb_ip7__T_5_mask = 1'h0;
  assign queue_bits_wb_ip7__T_5_en = 1'h0;
  assign queue_bits_wb_ip7__T_6_data = 1'h0;
  assign queue_bits_wb_ip7__T_6_addr = 6'h1;
  assign queue_bits_wb_ip7__T_6_mask = 1'h0;
  assign queue_bits_wb_ip7__T_6_en = 1'h0;
  assign queue_bits_wb_ip7__T_7_data = 1'h0;
  assign queue_bits_wb_ip7__T_7_addr = 6'h2;
  assign queue_bits_wb_ip7__T_7_mask = 1'h0;
  assign queue_bits_wb_ip7__T_7_en = 1'h0;
  assign queue_bits_wb_ip7__T_8_data = 1'h0;
  assign queue_bits_wb_ip7__T_8_addr = 6'h3;
  assign queue_bits_wb_ip7__T_8_mask = 1'h0;
  assign queue_bits_wb_ip7__T_8_en = 1'h0;
  assign queue_bits_wb_ip7__T_9_data = 1'h0;
  assign queue_bits_wb_ip7__T_9_addr = 6'h4;
  assign queue_bits_wb_ip7__T_9_mask = 1'h0;
  assign queue_bits_wb_ip7__T_9_en = 1'h0;
  assign queue_bits_wb_ip7__T_10_data = 1'h0;
  assign queue_bits_wb_ip7__T_10_addr = 6'h5;
  assign queue_bits_wb_ip7__T_10_mask = 1'h0;
  assign queue_bits_wb_ip7__T_10_en = 1'h0;
  assign queue_bits_wb_ip7__T_11_data = 1'h0;
  assign queue_bits_wb_ip7__T_11_addr = 6'h6;
  assign queue_bits_wb_ip7__T_11_mask = 1'h0;
  assign queue_bits_wb_ip7__T_11_en = 1'h0;
  assign queue_bits_wb_ip7__T_12_data = 1'h0;
  assign queue_bits_wb_ip7__T_12_addr = 6'h7;
  assign queue_bits_wb_ip7__T_12_mask = 1'h0;
  assign queue_bits_wb_ip7__T_12_en = 1'h0;
  assign queue_bits_wb_ip7__T_13_data = 1'h0;
  assign queue_bits_wb_ip7__T_13_addr = 6'h8;
  assign queue_bits_wb_ip7__T_13_mask = 1'h0;
  assign queue_bits_wb_ip7__T_13_en = 1'h0;
  assign queue_bits_wb_ip7__T_14_data = 1'h0;
  assign queue_bits_wb_ip7__T_14_addr = 6'h9;
  assign queue_bits_wb_ip7__T_14_mask = 1'h0;
  assign queue_bits_wb_ip7__T_14_en = 1'h0;
  assign queue_bits_wb_ip7__T_15_data = 1'h0;
  assign queue_bits_wb_ip7__T_15_addr = 6'ha;
  assign queue_bits_wb_ip7__T_15_mask = 1'h0;
  assign queue_bits_wb_ip7__T_15_en = 1'h0;
  assign queue_bits_wb_ip7__T_16_data = 1'h0;
  assign queue_bits_wb_ip7__T_16_addr = 6'hb;
  assign queue_bits_wb_ip7__T_16_mask = 1'h0;
  assign queue_bits_wb_ip7__T_16_en = 1'h0;
  assign queue_bits_wb_ip7__T_17_data = 1'h0;
  assign queue_bits_wb_ip7__T_17_addr = 6'hc;
  assign queue_bits_wb_ip7__T_17_mask = 1'h0;
  assign queue_bits_wb_ip7__T_17_en = 1'h0;
  assign queue_bits_wb_ip7__T_18_data = 1'h0;
  assign queue_bits_wb_ip7__T_18_addr = 6'hd;
  assign queue_bits_wb_ip7__T_18_mask = 1'h0;
  assign queue_bits_wb_ip7__T_18_en = 1'h0;
  assign queue_bits_wb_ip7__T_19_data = 1'h0;
  assign queue_bits_wb_ip7__T_19_addr = 6'he;
  assign queue_bits_wb_ip7__T_19_mask = 1'h0;
  assign queue_bits_wb_ip7__T_19_en = 1'h0;
  assign queue_bits_wb_ip7__T_20_data = 1'h0;
  assign queue_bits_wb_ip7__T_20_addr = 6'hf;
  assign queue_bits_wb_ip7__T_20_mask = 1'h0;
  assign queue_bits_wb_ip7__T_20_en = 1'h0;
  assign queue_bits_wb_ip7__T_21_data = 1'h0;
  assign queue_bits_wb_ip7__T_21_addr = 6'h10;
  assign queue_bits_wb_ip7__T_21_mask = 1'h0;
  assign queue_bits_wb_ip7__T_21_en = 1'h0;
  assign queue_bits_wb_ip7__T_22_data = 1'h0;
  assign queue_bits_wb_ip7__T_22_addr = 6'h11;
  assign queue_bits_wb_ip7__T_22_mask = 1'h0;
  assign queue_bits_wb_ip7__T_22_en = 1'h0;
  assign queue_bits_wb_ip7__T_23_data = 1'h0;
  assign queue_bits_wb_ip7__T_23_addr = 6'h12;
  assign queue_bits_wb_ip7__T_23_mask = 1'h0;
  assign queue_bits_wb_ip7__T_23_en = 1'h0;
  assign queue_bits_wb_ip7__T_24_data = 1'h0;
  assign queue_bits_wb_ip7__T_24_addr = 6'h13;
  assign queue_bits_wb_ip7__T_24_mask = 1'h0;
  assign queue_bits_wb_ip7__T_24_en = 1'h0;
  assign queue_bits_wb_ip7__T_25_data = 1'h0;
  assign queue_bits_wb_ip7__T_25_addr = 6'h14;
  assign queue_bits_wb_ip7__T_25_mask = 1'h0;
  assign queue_bits_wb_ip7__T_25_en = 1'h0;
  assign queue_bits_wb_ip7__T_26_data = 1'h0;
  assign queue_bits_wb_ip7__T_26_addr = 6'h15;
  assign queue_bits_wb_ip7__T_26_mask = 1'h0;
  assign queue_bits_wb_ip7__T_26_en = 1'h0;
  assign queue_bits_wb_ip7__T_27_data = 1'h0;
  assign queue_bits_wb_ip7__T_27_addr = 6'h16;
  assign queue_bits_wb_ip7__T_27_mask = 1'h0;
  assign queue_bits_wb_ip7__T_27_en = 1'h0;
  assign queue_bits_wb_ip7__T_28_data = 1'h0;
  assign queue_bits_wb_ip7__T_28_addr = 6'h17;
  assign queue_bits_wb_ip7__T_28_mask = 1'h0;
  assign queue_bits_wb_ip7__T_28_en = 1'h0;
  assign queue_bits_wb_ip7__T_29_data = 1'h0;
  assign queue_bits_wb_ip7__T_29_addr = 6'h18;
  assign queue_bits_wb_ip7__T_29_mask = 1'h0;
  assign queue_bits_wb_ip7__T_29_en = 1'h0;
  assign queue_bits_wb_ip7__T_30_data = 1'h0;
  assign queue_bits_wb_ip7__T_30_addr = 6'h19;
  assign queue_bits_wb_ip7__T_30_mask = 1'h0;
  assign queue_bits_wb_ip7__T_30_en = 1'h0;
  assign queue_bits_wb_ip7__T_31_data = 1'h0;
  assign queue_bits_wb_ip7__T_31_addr = 6'h1a;
  assign queue_bits_wb_ip7__T_31_mask = 1'h0;
  assign queue_bits_wb_ip7__T_31_en = 1'h0;
  assign queue_bits_wb_ip7__T_32_data = 1'h0;
  assign queue_bits_wb_ip7__T_32_addr = 6'h1b;
  assign queue_bits_wb_ip7__T_32_mask = 1'h0;
  assign queue_bits_wb_ip7__T_32_en = 1'h0;
  assign queue_bits_wb_ip7__T_33_data = 1'h0;
  assign queue_bits_wb_ip7__T_33_addr = 6'h1c;
  assign queue_bits_wb_ip7__T_33_mask = 1'h0;
  assign queue_bits_wb_ip7__T_33_en = 1'h0;
  assign queue_bits_wb_ip7__T_34_data = 1'h0;
  assign queue_bits_wb_ip7__T_34_addr = 6'h1d;
  assign queue_bits_wb_ip7__T_34_mask = 1'h0;
  assign queue_bits_wb_ip7__T_34_en = 1'h0;
  assign queue_bits_wb_ip7__T_35_data = 1'h0;
  assign queue_bits_wb_ip7__T_35_addr = 6'h1e;
  assign queue_bits_wb_ip7__T_35_mask = 1'h0;
  assign queue_bits_wb_ip7__T_35_en = 1'h0;
  assign queue_bits_wb_ip7__T_36_data = 1'h0;
  assign queue_bits_wb_ip7__T_36_addr = 6'h1f;
  assign queue_bits_wb_ip7__T_36_mask = 1'h0;
  assign queue_bits_wb_ip7__T_36_en = 1'h0;
  assign queue_bits_wb_ip7__T_37_data = 1'h0;
  assign queue_bits_wb_ip7__T_37_addr = 6'h20;
  assign queue_bits_wb_ip7__T_37_mask = 1'h0;
  assign queue_bits_wb_ip7__T_37_en = 1'h0;
  assign queue_bits_wb_ip7__T_38_data = 1'h0;
  assign queue_bits_wb_ip7__T_38_addr = 6'h21;
  assign queue_bits_wb_ip7__T_38_mask = 1'h0;
  assign queue_bits_wb_ip7__T_38_en = 1'h0;
  assign queue_bits_wb_ip7__T_39_data = 1'h0;
  assign queue_bits_wb_ip7__T_39_addr = 6'h22;
  assign queue_bits_wb_ip7__T_39_mask = 1'h0;
  assign queue_bits_wb_ip7__T_39_en = 1'h0;
  assign queue_bits_wb_ip7__T_40_data = 1'h0;
  assign queue_bits_wb_ip7__T_40_addr = 6'h23;
  assign queue_bits_wb_ip7__T_40_mask = 1'h0;
  assign queue_bits_wb_ip7__T_40_en = 1'h0;
  assign queue_bits_wb_ip7__T_41_data = 1'h0;
  assign queue_bits_wb_ip7__T_41_addr = 6'h24;
  assign queue_bits_wb_ip7__T_41_mask = 1'h0;
  assign queue_bits_wb_ip7__T_41_en = 1'h0;
  assign queue_bits_wb_ip7__T_42_data = 1'h0;
  assign queue_bits_wb_ip7__T_42_addr = 6'h25;
  assign queue_bits_wb_ip7__T_42_mask = 1'h0;
  assign queue_bits_wb_ip7__T_42_en = 1'h0;
  assign queue_bits_wb_ip7__T_43_data = 1'h0;
  assign queue_bits_wb_ip7__T_43_addr = 6'h26;
  assign queue_bits_wb_ip7__T_43_mask = 1'h0;
  assign queue_bits_wb_ip7__T_43_en = 1'h0;
  assign queue_bits_wb_ip7__T_44_data = 1'h0;
  assign queue_bits_wb_ip7__T_44_addr = 6'h27;
  assign queue_bits_wb_ip7__T_44_mask = 1'h0;
  assign queue_bits_wb_ip7__T_44_en = 1'h0;
  assign queue_bits_wb_ip7__T_45_data = 1'h0;
  assign queue_bits_wb_ip7__T_45_addr = 6'h28;
  assign queue_bits_wb_ip7__T_45_mask = 1'h0;
  assign queue_bits_wb_ip7__T_45_en = 1'h0;
  assign queue_bits_wb_ip7__T_46_data = 1'h0;
  assign queue_bits_wb_ip7__T_46_addr = 6'h29;
  assign queue_bits_wb_ip7__T_46_mask = 1'h0;
  assign queue_bits_wb_ip7__T_46_en = 1'h0;
  assign queue_bits_wb_ip7__T_47_data = 1'h0;
  assign queue_bits_wb_ip7__T_47_addr = 6'h2a;
  assign queue_bits_wb_ip7__T_47_mask = 1'h0;
  assign queue_bits_wb_ip7__T_47_en = 1'h0;
  assign queue_bits_wb_ip7__T_48_data = 1'h0;
  assign queue_bits_wb_ip7__T_48_addr = 6'h2b;
  assign queue_bits_wb_ip7__T_48_mask = 1'h0;
  assign queue_bits_wb_ip7__T_48_en = 1'h0;
  assign queue_bits_wb_ip7__T_49_data = 1'h0;
  assign queue_bits_wb_ip7__T_49_addr = 6'h2c;
  assign queue_bits_wb_ip7__T_49_mask = 1'h0;
  assign queue_bits_wb_ip7__T_49_en = 1'h0;
  assign queue_bits_wb_ip7__T_50_data = 1'h0;
  assign queue_bits_wb_ip7__T_50_addr = 6'h2d;
  assign queue_bits_wb_ip7__T_50_mask = 1'h0;
  assign queue_bits_wb_ip7__T_50_en = 1'h0;
  assign queue_bits_wb_ip7__T_51_data = 1'h0;
  assign queue_bits_wb_ip7__T_51_addr = 6'h2e;
  assign queue_bits_wb_ip7__T_51_mask = 1'h0;
  assign queue_bits_wb_ip7__T_51_en = 1'h0;
  assign queue_bits_wb_ip7__T_52_data = 1'h0;
  assign queue_bits_wb_ip7__T_52_addr = 6'h2f;
  assign queue_bits_wb_ip7__T_52_mask = 1'h0;
  assign queue_bits_wb_ip7__T_52_en = 1'h0;
  assign queue_bits_wb_ip7__T_53_data = 1'h0;
  assign queue_bits_wb_ip7__T_53_addr = 6'h30;
  assign queue_bits_wb_ip7__T_53_mask = 1'h0;
  assign queue_bits_wb_ip7__T_53_en = 1'h0;
  assign queue_bits_wb_ip7__T_54_data = 1'h0;
  assign queue_bits_wb_ip7__T_54_addr = 6'h31;
  assign queue_bits_wb_ip7__T_54_mask = 1'h0;
  assign queue_bits_wb_ip7__T_54_en = 1'h0;
  assign queue_bits_wb_ip7__T_55_data = 1'h0;
  assign queue_bits_wb_ip7__T_55_addr = 6'h32;
  assign queue_bits_wb_ip7__T_55_mask = 1'h0;
  assign queue_bits_wb_ip7__T_55_en = 1'h0;
  assign queue_bits_wb_ip7__T_56_data = 1'h0;
  assign queue_bits_wb_ip7__T_56_addr = 6'h33;
  assign queue_bits_wb_ip7__T_56_mask = 1'h0;
  assign queue_bits_wb_ip7__T_56_en = 1'h0;
  assign queue_bits_wb_ip7__T_57_data = 1'h0;
  assign queue_bits_wb_ip7__T_57_addr = 6'h34;
  assign queue_bits_wb_ip7__T_57_mask = 1'h0;
  assign queue_bits_wb_ip7__T_57_en = 1'h0;
  assign queue_bits_wb_ip7__T_58_data = 1'h0;
  assign queue_bits_wb_ip7__T_58_addr = 6'h35;
  assign queue_bits_wb_ip7__T_58_mask = 1'h0;
  assign queue_bits_wb_ip7__T_58_en = 1'h0;
  assign queue_bits_wb_ip7__T_59_data = 1'h0;
  assign queue_bits_wb_ip7__T_59_addr = 6'h36;
  assign queue_bits_wb_ip7__T_59_mask = 1'h0;
  assign queue_bits_wb_ip7__T_59_en = 1'h0;
  assign queue_bits_wb_ip7__T_60_data = 1'h0;
  assign queue_bits_wb_ip7__T_60_addr = 6'h37;
  assign queue_bits_wb_ip7__T_60_mask = 1'h0;
  assign queue_bits_wb_ip7__T_60_en = 1'h0;
  assign queue_bits_wb_ip7__T_61_data = 1'h0;
  assign queue_bits_wb_ip7__T_61_addr = 6'h38;
  assign queue_bits_wb_ip7__T_61_mask = 1'h0;
  assign queue_bits_wb_ip7__T_61_en = 1'h0;
  assign queue_bits_wb_ip7__T_62_data = 1'h0;
  assign queue_bits_wb_ip7__T_62_addr = 6'h39;
  assign queue_bits_wb_ip7__T_62_mask = 1'h0;
  assign queue_bits_wb_ip7__T_62_en = 1'h0;
  assign queue_bits_wb_ip7__T_63_data = 1'h0;
  assign queue_bits_wb_ip7__T_63_addr = 6'h3a;
  assign queue_bits_wb_ip7__T_63_mask = 1'h0;
  assign queue_bits_wb_ip7__T_63_en = 1'h0;
  assign queue_bits_wb_ip7__T_64_data = 1'h0;
  assign queue_bits_wb_ip7__T_64_addr = 6'h3b;
  assign queue_bits_wb_ip7__T_64_mask = 1'h0;
  assign queue_bits_wb_ip7__T_64_en = 1'h0;
  assign queue_bits_wb_ip7__T_65_data = 1'h0;
  assign queue_bits_wb_ip7__T_65_addr = 6'h3c;
  assign queue_bits_wb_ip7__T_65_mask = 1'h0;
  assign queue_bits_wb_ip7__T_65_en = 1'h0;
  assign queue_bits_wb_ip7__T_66_data = 1'h0;
  assign queue_bits_wb_ip7__T_66_addr = 6'h3d;
  assign queue_bits_wb_ip7__T_66_mask = 1'h0;
  assign queue_bits_wb_ip7__T_66_en = 1'h0;
  assign queue_bits_wb_ip7__T_67_data = 1'h0;
  assign queue_bits_wb_ip7__T_67_addr = 6'h3e;
  assign queue_bits_wb_ip7__T_67_mask = 1'h0;
  assign queue_bits_wb_ip7__T_67_en = 1'h0;
  assign queue_bits_wb_ip7__T_68_data = 1'h0;
  assign queue_bits_wb_ip7__T_68_addr = 6'h3f;
  assign queue_bits_wb_ip7__T_68_mask = 1'h0;
  assign queue_bits_wb_ip7__T_68_en = 1'h0;
  assign queue_bits_wb_ip7__T_70_data = 1'h0;
  assign queue_bits_wb_ip7__T_70_addr = 6'h0;
  assign queue_bits_wb_ip7__T_70_mask = 1'h0;
  assign queue_bits_wb_ip7__T_70_en = reset;
  assign queue_bits_wb_ip7__T_71_data = 1'h0;
  assign queue_bits_wb_ip7__T_71_addr = 6'h1;
  assign queue_bits_wb_ip7__T_71_mask = 1'h0;
  assign queue_bits_wb_ip7__T_71_en = reset;
  assign queue_bits_wb_ip7__T_72_data = 1'h0;
  assign queue_bits_wb_ip7__T_72_addr = 6'h2;
  assign queue_bits_wb_ip7__T_72_mask = 1'h0;
  assign queue_bits_wb_ip7__T_72_en = reset;
  assign queue_bits_wb_ip7__T_73_data = 1'h0;
  assign queue_bits_wb_ip7__T_73_addr = 6'h3;
  assign queue_bits_wb_ip7__T_73_mask = 1'h0;
  assign queue_bits_wb_ip7__T_73_en = reset;
  assign queue_bits_wb_ip7__T_74_data = 1'h0;
  assign queue_bits_wb_ip7__T_74_addr = 6'h4;
  assign queue_bits_wb_ip7__T_74_mask = 1'h0;
  assign queue_bits_wb_ip7__T_74_en = reset;
  assign queue_bits_wb_ip7__T_75_data = 1'h0;
  assign queue_bits_wb_ip7__T_75_addr = 6'h5;
  assign queue_bits_wb_ip7__T_75_mask = 1'h0;
  assign queue_bits_wb_ip7__T_75_en = reset;
  assign queue_bits_wb_ip7__T_76_data = 1'h0;
  assign queue_bits_wb_ip7__T_76_addr = 6'h6;
  assign queue_bits_wb_ip7__T_76_mask = 1'h0;
  assign queue_bits_wb_ip7__T_76_en = reset;
  assign queue_bits_wb_ip7__T_77_data = 1'h0;
  assign queue_bits_wb_ip7__T_77_addr = 6'h7;
  assign queue_bits_wb_ip7__T_77_mask = 1'h0;
  assign queue_bits_wb_ip7__T_77_en = reset;
  assign queue_bits_wb_ip7__T_78_data = 1'h0;
  assign queue_bits_wb_ip7__T_78_addr = 6'h8;
  assign queue_bits_wb_ip7__T_78_mask = 1'h0;
  assign queue_bits_wb_ip7__T_78_en = reset;
  assign queue_bits_wb_ip7__T_79_data = 1'h0;
  assign queue_bits_wb_ip7__T_79_addr = 6'h9;
  assign queue_bits_wb_ip7__T_79_mask = 1'h0;
  assign queue_bits_wb_ip7__T_79_en = reset;
  assign queue_bits_wb_ip7__T_80_data = 1'h0;
  assign queue_bits_wb_ip7__T_80_addr = 6'ha;
  assign queue_bits_wb_ip7__T_80_mask = 1'h0;
  assign queue_bits_wb_ip7__T_80_en = reset;
  assign queue_bits_wb_ip7__T_81_data = 1'h0;
  assign queue_bits_wb_ip7__T_81_addr = 6'hb;
  assign queue_bits_wb_ip7__T_81_mask = 1'h0;
  assign queue_bits_wb_ip7__T_81_en = reset;
  assign queue_bits_wb_ip7__T_82_data = 1'h0;
  assign queue_bits_wb_ip7__T_82_addr = 6'hc;
  assign queue_bits_wb_ip7__T_82_mask = 1'h0;
  assign queue_bits_wb_ip7__T_82_en = reset;
  assign queue_bits_wb_ip7__T_83_data = 1'h0;
  assign queue_bits_wb_ip7__T_83_addr = 6'hd;
  assign queue_bits_wb_ip7__T_83_mask = 1'h0;
  assign queue_bits_wb_ip7__T_83_en = reset;
  assign queue_bits_wb_ip7__T_84_data = 1'h0;
  assign queue_bits_wb_ip7__T_84_addr = 6'he;
  assign queue_bits_wb_ip7__T_84_mask = 1'h0;
  assign queue_bits_wb_ip7__T_84_en = reset;
  assign queue_bits_wb_ip7__T_85_data = 1'h0;
  assign queue_bits_wb_ip7__T_85_addr = 6'hf;
  assign queue_bits_wb_ip7__T_85_mask = 1'h0;
  assign queue_bits_wb_ip7__T_85_en = reset;
  assign queue_bits_wb_ip7__T_86_data = 1'h0;
  assign queue_bits_wb_ip7__T_86_addr = 6'h10;
  assign queue_bits_wb_ip7__T_86_mask = 1'h0;
  assign queue_bits_wb_ip7__T_86_en = reset;
  assign queue_bits_wb_ip7__T_87_data = 1'h0;
  assign queue_bits_wb_ip7__T_87_addr = 6'h11;
  assign queue_bits_wb_ip7__T_87_mask = 1'h0;
  assign queue_bits_wb_ip7__T_87_en = reset;
  assign queue_bits_wb_ip7__T_88_data = 1'h0;
  assign queue_bits_wb_ip7__T_88_addr = 6'h12;
  assign queue_bits_wb_ip7__T_88_mask = 1'h0;
  assign queue_bits_wb_ip7__T_88_en = reset;
  assign queue_bits_wb_ip7__T_89_data = 1'h0;
  assign queue_bits_wb_ip7__T_89_addr = 6'h13;
  assign queue_bits_wb_ip7__T_89_mask = 1'h0;
  assign queue_bits_wb_ip7__T_89_en = reset;
  assign queue_bits_wb_ip7__T_90_data = 1'h0;
  assign queue_bits_wb_ip7__T_90_addr = 6'h14;
  assign queue_bits_wb_ip7__T_90_mask = 1'h0;
  assign queue_bits_wb_ip7__T_90_en = reset;
  assign queue_bits_wb_ip7__T_91_data = 1'h0;
  assign queue_bits_wb_ip7__T_91_addr = 6'h15;
  assign queue_bits_wb_ip7__T_91_mask = 1'h0;
  assign queue_bits_wb_ip7__T_91_en = reset;
  assign queue_bits_wb_ip7__T_92_data = 1'h0;
  assign queue_bits_wb_ip7__T_92_addr = 6'h16;
  assign queue_bits_wb_ip7__T_92_mask = 1'h0;
  assign queue_bits_wb_ip7__T_92_en = reset;
  assign queue_bits_wb_ip7__T_93_data = 1'h0;
  assign queue_bits_wb_ip7__T_93_addr = 6'h17;
  assign queue_bits_wb_ip7__T_93_mask = 1'h0;
  assign queue_bits_wb_ip7__T_93_en = reset;
  assign queue_bits_wb_ip7__T_94_data = 1'h0;
  assign queue_bits_wb_ip7__T_94_addr = 6'h18;
  assign queue_bits_wb_ip7__T_94_mask = 1'h0;
  assign queue_bits_wb_ip7__T_94_en = reset;
  assign queue_bits_wb_ip7__T_95_data = 1'h0;
  assign queue_bits_wb_ip7__T_95_addr = 6'h19;
  assign queue_bits_wb_ip7__T_95_mask = 1'h0;
  assign queue_bits_wb_ip7__T_95_en = reset;
  assign queue_bits_wb_ip7__T_96_data = 1'h0;
  assign queue_bits_wb_ip7__T_96_addr = 6'h1a;
  assign queue_bits_wb_ip7__T_96_mask = 1'h0;
  assign queue_bits_wb_ip7__T_96_en = reset;
  assign queue_bits_wb_ip7__T_97_data = 1'h0;
  assign queue_bits_wb_ip7__T_97_addr = 6'h1b;
  assign queue_bits_wb_ip7__T_97_mask = 1'h0;
  assign queue_bits_wb_ip7__T_97_en = reset;
  assign queue_bits_wb_ip7__T_98_data = 1'h0;
  assign queue_bits_wb_ip7__T_98_addr = 6'h1c;
  assign queue_bits_wb_ip7__T_98_mask = 1'h0;
  assign queue_bits_wb_ip7__T_98_en = reset;
  assign queue_bits_wb_ip7__T_99_data = 1'h0;
  assign queue_bits_wb_ip7__T_99_addr = 6'h1d;
  assign queue_bits_wb_ip7__T_99_mask = 1'h0;
  assign queue_bits_wb_ip7__T_99_en = reset;
  assign queue_bits_wb_ip7__T_100_data = 1'h0;
  assign queue_bits_wb_ip7__T_100_addr = 6'h1e;
  assign queue_bits_wb_ip7__T_100_mask = 1'h0;
  assign queue_bits_wb_ip7__T_100_en = reset;
  assign queue_bits_wb_ip7__T_101_data = 1'h0;
  assign queue_bits_wb_ip7__T_101_addr = 6'h1f;
  assign queue_bits_wb_ip7__T_101_mask = 1'h0;
  assign queue_bits_wb_ip7__T_101_en = reset;
  assign queue_bits_wb_ip7__T_102_data = 1'h0;
  assign queue_bits_wb_ip7__T_102_addr = 6'h20;
  assign queue_bits_wb_ip7__T_102_mask = 1'h0;
  assign queue_bits_wb_ip7__T_102_en = reset;
  assign queue_bits_wb_ip7__T_103_data = 1'h0;
  assign queue_bits_wb_ip7__T_103_addr = 6'h21;
  assign queue_bits_wb_ip7__T_103_mask = 1'h0;
  assign queue_bits_wb_ip7__T_103_en = reset;
  assign queue_bits_wb_ip7__T_104_data = 1'h0;
  assign queue_bits_wb_ip7__T_104_addr = 6'h22;
  assign queue_bits_wb_ip7__T_104_mask = 1'h0;
  assign queue_bits_wb_ip7__T_104_en = reset;
  assign queue_bits_wb_ip7__T_105_data = 1'h0;
  assign queue_bits_wb_ip7__T_105_addr = 6'h23;
  assign queue_bits_wb_ip7__T_105_mask = 1'h0;
  assign queue_bits_wb_ip7__T_105_en = reset;
  assign queue_bits_wb_ip7__T_106_data = 1'h0;
  assign queue_bits_wb_ip7__T_106_addr = 6'h24;
  assign queue_bits_wb_ip7__T_106_mask = 1'h0;
  assign queue_bits_wb_ip7__T_106_en = reset;
  assign queue_bits_wb_ip7__T_107_data = 1'h0;
  assign queue_bits_wb_ip7__T_107_addr = 6'h25;
  assign queue_bits_wb_ip7__T_107_mask = 1'h0;
  assign queue_bits_wb_ip7__T_107_en = reset;
  assign queue_bits_wb_ip7__T_108_data = 1'h0;
  assign queue_bits_wb_ip7__T_108_addr = 6'h26;
  assign queue_bits_wb_ip7__T_108_mask = 1'h0;
  assign queue_bits_wb_ip7__T_108_en = reset;
  assign queue_bits_wb_ip7__T_109_data = 1'h0;
  assign queue_bits_wb_ip7__T_109_addr = 6'h27;
  assign queue_bits_wb_ip7__T_109_mask = 1'h0;
  assign queue_bits_wb_ip7__T_109_en = reset;
  assign queue_bits_wb_ip7__T_110_data = 1'h0;
  assign queue_bits_wb_ip7__T_110_addr = 6'h28;
  assign queue_bits_wb_ip7__T_110_mask = 1'h0;
  assign queue_bits_wb_ip7__T_110_en = reset;
  assign queue_bits_wb_ip7__T_111_data = 1'h0;
  assign queue_bits_wb_ip7__T_111_addr = 6'h29;
  assign queue_bits_wb_ip7__T_111_mask = 1'h0;
  assign queue_bits_wb_ip7__T_111_en = reset;
  assign queue_bits_wb_ip7__T_112_data = 1'h0;
  assign queue_bits_wb_ip7__T_112_addr = 6'h2a;
  assign queue_bits_wb_ip7__T_112_mask = 1'h0;
  assign queue_bits_wb_ip7__T_112_en = reset;
  assign queue_bits_wb_ip7__T_113_data = 1'h0;
  assign queue_bits_wb_ip7__T_113_addr = 6'h2b;
  assign queue_bits_wb_ip7__T_113_mask = 1'h0;
  assign queue_bits_wb_ip7__T_113_en = reset;
  assign queue_bits_wb_ip7__T_114_data = 1'h0;
  assign queue_bits_wb_ip7__T_114_addr = 6'h2c;
  assign queue_bits_wb_ip7__T_114_mask = 1'h0;
  assign queue_bits_wb_ip7__T_114_en = reset;
  assign queue_bits_wb_ip7__T_115_data = 1'h0;
  assign queue_bits_wb_ip7__T_115_addr = 6'h2d;
  assign queue_bits_wb_ip7__T_115_mask = 1'h0;
  assign queue_bits_wb_ip7__T_115_en = reset;
  assign queue_bits_wb_ip7__T_116_data = 1'h0;
  assign queue_bits_wb_ip7__T_116_addr = 6'h2e;
  assign queue_bits_wb_ip7__T_116_mask = 1'h0;
  assign queue_bits_wb_ip7__T_116_en = reset;
  assign queue_bits_wb_ip7__T_117_data = 1'h0;
  assign queue_bits_wb_ip7__T_117_addr = 6'h2f;
  assign queue_bits_wb_ip7__T_117_mask = 1'h0;
  assign queue_bits_wb_ip7__T_117_en = reset;
  assign queue_bits_wb_ip7__T_118_data = 1'h0;
  assign queue_bits_wb_ip7__T_118_addr = 6'h30;
  assign queue_bits_wb_ip7__T_118_mask = 1'h0;
  assign queue_bits_wb_ip7__T_118_en = reset;
  assign queue_bits_wb_ip7__T_119_data = 1'h0;
  assign queue_bits_wb_ip7__T_119_addr = 6'h31;
  assign queue_bits_wb_ip7__T_119_mask = 1'h0;
  assign queue_bits_wb_ip7__T_119_en = reset;
  assign queue_bits_wb_ip7__T_120_data = 1'h0;
  assign queue_bits_wb_ip7__T_120_addr = 6'h32;
  assign queue_bits_wb_ip7__T_120_mask = 1'h0;
  assign queue_bits_wb_ip7__T_120_en = reset;
  assign queue_bits_wb_ip7__T_121_data = 1'h0;
  assign queue_bits_wb_ip7__T_121_addr = 6'h33;
  assign queue_bits_wb_ip7__T_121_mask = 1'h0;
  assign queue_bits_wb_ip7__T_121_en = reset;
  assign queue_bits_wb_ip7__T_122_data = 1'h0;
  assign queue_bits_wb_ip7__T_122_addr = 6'h34;
  assign queue_bits_wb_ip7__T_122_mask = 1'h0;
  assign queue_bits_wb_ip7__T_122_en = reset;
  assign queue_bits_wb_ip7__T_123_data = 1'h0;
  assign queue_bits_wb_ip7__T_123_addr = 6'h35;
  assign queue_bits_wb_ip7__T_123_mask = 1'h0;
  assign queue_bits_wb_ip7__T_123_en = reset;
  assign queue_bits_wb_ip7__T_124_data = 1'h0;
  assign queue_bits_wb_ip7__T_124_addr = 6'h36;
  assign queue_bits_wb_ip7__T_124_mask = 1'h0;
  assign queue_bits_wb_ip7__T_124_en = reset;
  assign queue_bits_wb_ip7__T_125_data = 1'h0;
  assign queue_bits_wb_ip7__T_125_addr = 6'h37;
  assign queue_bits_wb_ip7__T_125_mask = 1'h0;
  assign queue_bits_wb_ip7__T_125_en = reset;
  assign queue_bits_wb_ip7__T_126_data = 1'h0;
  assign queue_bits_wb_ip7__T_126_addr = 6'h38;
  assign queue_bits_wb_ip7__T_126_mask = 1'h0;
  assign queue_bits_wb_ip7__T_126_en = reset;
  assign queue_bits_wb_ip7__T_127_data = 1'h0;
  assign queue_bits_wb_ip7__T_127_addr = 6'h39;
  assign queue_bits_wb_ip7__T_127_mask = 1'h0;
  assign queue_bits_wb_ip7__T_127_en = reset;
  assign queue_bits_wb_ip7__T_128_data = 1'h0;
  assign queue_bits_wb_ip7__T_128_addr = 6'h3a;
  assign queue_bits_wb_ip7__T_128_mask = 1'h0;
  assign queue_bits_wb_ip7__T_128_en = reset;
  assign queue_bits_wb_ip7__T_129_data = 1'h0;
  assign queue_bits_wb_ip7__T_129_addr = 6'h3b;
  assign queue_bits_wb_ip7__T_129_mask = 1'h0;
  assign queue_bits_wb_ip7__T_129_en = reset;
  assign queue_bits_wb_ip7__T_130_data = 1'h0;
  assign queue_bits_wb_ip7__T_130_addr = 6'h3c;
  assign queue_bits_wb_ip7__T_130_mask = 1'h0;
  assign queue_bits_wb_ip7__T_130_en = reset;
  assign queue_bits_wb_ip7__T_131_data = 1'h0;
  assign queue_bits_wb_ip7__T_131_addr = 6'h3d;
  assign queue_bits_wb_ip7__T_131_mask = 1'h0;
  assign queue_bits_wb_ip7__T_131_en = reset;
  assign queue_bits_wb_ip7__T_132_data = 1'h0;
  assign queue_bits_wb_ip7__T_132_addr = 6'h3e;
  assign queue_bits_wb_ip7__T_132_mask = 1'h0;
  assign queue_bits_wb_ip7__T_132_en = reset;
  assign queue_bits_wb_ip7__T_133_data = 1'h0;
  assign queue_bits_wb_ip7__T_133_addr = 6'h3f;
  assign queue_bits_wb_ip7__T_133_mask = 1'h0;
  assign queue_bits_wb_ip7__T_133_en = reset;
  assign queue_bits_wb_ip7_q_head_w_data = 1'h0;
  assign queue_bits_wb_ip7_q_head_w_addr = head;
  assign queue_bits_wb_ip7_q_head_w_mask = 1'h0;
  assign queue_bits_wb_ip7_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_is_ds_q_head_r_addr = head;
  assign queue_bits_wb_is_ds_q_head_r_data = queue_bits_wb_is_ds[queue_bits_wb_is_ds_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_is_ds__T_3_data = io_enq_0_bits_data_wb_is_ds;
  assign queue_bits_wb_is_ds__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_is_ds__T_3_mask = 1'h1;
  assign queue_bits_wb_is_ds__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_is_ds__T_4_data = io_enq_1_bits_data_wb_is_ds;
  assign queue_bits_wb_is_ds__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_is_ds__T_4_mask = 1'h1;
  assign queue_bits_wb_is_ds__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_is_ds__T_5_data = 1'h0;
  assign queue_bits_wb_is_ds__T_5_addr = 6'h0;
  assign queue_bits_wb_is_ds__T_5_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_5_en = 1'h0;
  assign queue_bits_wb_is_ds__T_6_data = 1'h0;
  assign queue_bits_wb_is_ds__T_6_addr = 6'h1;
  assign queue_bits_wb_is_ds__T_6_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_6_en = 1'h0;
  assign queue_bits_wb_is_ds__T_7_data = 1'h0;
  assign queue_bits_wb_is_ds__T_7_addr = 6'h2;
  assign queue_bits_wb_is_ds__T_7_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_7_en = 1'h0;
  assign queue_bits_wb_is_ds__T_8_data = 1'h0;
  assign queue_bits_wb_is_ds__T_8_addr = 6'h3;
  assign queue_bits_wb_is_ds__T_8_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_8_en = 1'h0;
  assign queue_bits_wb_is_ds__T_9_data = 1'h0;
  assign queue_bits_wb_is_ds__T_9_addr = 6'h4;
  assign queue_bits_wb_is_ds__T_9_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_9_en = 1'h0;
  assign queue_bits_wb_is_ds__T_10_data = 1'h0;
  assign queue_bits_wb_is_ds__T_10_addr = 6'h5;
  assign queue_bits_wb_is_ds__T_10_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_10_en = 1'h0;
  assign queue_bits_wb_is_ds__T_11_data = 1'h0;
  assign queue_bits_wb_is_ds__T_11_addr = 6'h6;
  assign queue_bits_wb_is_ds__T_11_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_11_en = 1'h0;
  assign queue_bits_wb_is_ds__T_12_data = 1'h0;
  assign queue_bits_wb_is_ds__T_12_addr = 6'h7;
  assign queue_bits_wb_is_ds__T_12_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_12_en = 1'h0;
  assign queue_bits_wb_is_ds__T_13_data = 1'h0;
  assign queue_bits_wb_is_ds__T_13_addr = 6'h8;
  assign queue_bits_wb_is_ds__T_13_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_13_en = 1'h0;
  assign queue_bits_wb_is_ds__T_14_data = 1'h0;
  assign queue_bits_wb_is_ds__T_14_addr = 6'h9;
  assign queue_bits_wb_is_ds__T_14_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_14_en = 1'h0;
  assign queue_bits_wb_is_ds__T_15_data = 1'h0;
  assign queue_bits_wb_is_ds__T_15_addr = 6'ha;
  assign queue_bits_wb_is_ds__T_15_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_15_en = 1'h0;
  assign queue_bits_wb_is_ds__T_16_data = 1'h0;
  assign queue_bits_wb_is_ds__T_16_addr = 6'hb;
  assign queue_bits_wb_is_ds__T_16_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_16_en = 1'h0;
  assign queue_bits_wb_is_ds__T_17_data = 1'h0;
  assign queue_bits_wb_is_ds__T_17_addr = 6'hc;
  assign queue_bits_wb_is_ds__T_17_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_17_en = 1'h0;
  assign queue_bits_wb_is_ds__T_18_data = 1'h0;
  assign queue_bits_wb_is_ds__T_18_addr = 6'hd;
  assign queue_bits_wb_is_ds__T_18_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_18_en = 1'h0;
  assign queue_bits_wb_is_ds__T_19_data = 1'h0;
  assign queue_bits_wb_is_ds__T_19_addr = 6'he;
  assign queue_bits_wb_is_ds__T_19_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_19_en = 1'h0;
  assign queue_bits_wb_is_ds__T_20_data = 1'h0;
  assign queue_bits_wb_is_ds__T_20_addr = 6'hf;
  assign queue_bits_wb_is_ds__T_20_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_20_en = 1'h0;
  assign queue_bits_wb_is_ds__T_21_data = 1'h0;
  assign queue_bits_wb_is_ds__T_21_addr = 6'h10;
  assign queue_bits_wb_is_ds__T_21_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_21_en = 1'h0;
  assign queue_bits_wb_is_ds__T_22_data = 1'h0;
  assign queue_bits_wb_is_ds__T_22_addr = 6'h11;
  assign queue_bits_wb_is_ds__T_22_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_22_en = 1'h0;
  assign queue_bits_wb_is_ds__T_23_data = 1'h0;
  assign queue_bits_wb_is_ds__T_23_addr = 6'h12;
  assign queue_bits_wb_is_ds__T_23_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_23_en = 1'h0;
  assign queue_bits_wb_is_ds__T_24_data = 1'h0;
  assign queue_bits_wb_is_ds__T_24_addr = 6'h13;
  assign queue_bits_wb_is_ds__T_24_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_24_en = 1'h0;
  assign queue_bits_wb_is_ds__T_25_data = 1'h0;
  assign queue_bits_wb_is_ds__T_25_addr = 6'h14;
  assign queue_bits_wb_is_ds__T_25_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_25_en = 1'h0;
  assign queue_bits_wb_is_ds__T_26_data = 1'h0;
  assign queue_bits_wb_is_ds__T_26_addr = 6'h15;
  assign queue_bits_wb_is_ds__T_26_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_26_en = 1'h0;
  assign queue_bits_wb_is_ds__T_27_data = 1'h0;
  assign queue_bits_wb_is_ds__T_27_addr = 6'h16;
  assign queue_bits_wb_is_ds__T_27_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_27_en = 1'h0;
  assign queue_bits_wb_is_ds__T_28_data = 1'h0;
  assign queue_bits_wb_is_ds__T_28_addr = 6'h17;
  assign queue_bits_wb_is_ds__T_28_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_28_en = 1'h0;
  assign queue_bits_wb_is_ds__T_29_data = 1'h0;
  assign queue_bits_wb_is_ds__T_29_addr = 6'h18;
  assign queue_bits_wb_is_ds__T_29_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_29_en = 1'h0;
  assign queue_bits_wb_is_ds__T_30_data = 1'h0;
  assign queue_bits_wb_is_ds__T_30_addr = 6'h19;
  assign queue_bits_wb_is_ds__T_30_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_30_en = 1'h0;
  assign queue_bits_wb_is_ds__T_31_data = 1'h0;
  assign queue_bits_wb_is_ds__T_31_addr = 6'h1a;
  assign queue_bits_wb_is_ds__T_31_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_31_en = 1'h0;
  assign queue_bits_wb_is_ds__T_32_data = 1'h0;
  assign queue_bits_wb_is_ds__T_32_addr = 6'h1b;
  assign queue_bits_wb_is_ds__T_32_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_32_en = 1'h0;
  assign queue_bits_wb_is_ds__T_33_data = 1'h0;
  assign queue_bits_wb_is_ds__T_33_addr = 6'h1c;
  assign queue_bits_wb_is_ds__T_33_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_33_en = 1'h0;
  assign queue_bits_wb_is_ds__T_34_data = 1'h0;
  assign queue_bits_wb_is_ds__T_34_addr = 6'h1d;
  assign queue_bits_wb_is_ds__T_34_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_34_en = 1'h0;
  assign queue_bits_wb_is_ds__T_35_data = 1'h0;
  assign queue_bits_wb_is_ds__T_35_addr = 6'h1e;
  assign queue_bits_wb_is_ds__T_35_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_35_en = 1'h0;
  assign queue_bits_wb_is_ds__T_36_data = 1'h0;
  assign queue_bits_wb_is_ds__T_36_addr = 6'h1f;
  assign queue_bits_wb_is_ds__T_36_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_36_en = 1'h0;
  assign queue_bits_wb_is_ds__T_37_data = 1'h0;
  assign queue_bits_wb_is_ds__T_37_addr = 6'h20;
  assign queue_bits_wb_is_ds__T_37_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_37_en = 1'h0;
  assign queue_bits_wb_is_ds__T_38_data = 1'h0;
  assign queue_bits_wb_is_ds__T_38_addr = 6'h21;
  assign queue_bits_wb_is_ds__T_38_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_38_en = 1'h0;
  assign queue_bits_wb_is_ds__T_39_data = 1'h0;
  assign queue_bits_wb_is_ds__T_39_addr = 6'h22;
  assign queue_bits_wb_is_ds__T_39_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_39_en = 1'h0;
  assign queue_bits_wb_is_ds__T_40_data = 1'h0;
  assign queue_bits_wb_is_ds__T_40_addr = 6'h23;
  assign queue_bits_wb_is_ds__T_40_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_40_en = 1'h0;
  assign queue_bits_wb_is_ds__T_41_data = 1'h0;
  assign queue_bits_wb_is_ds__T_41_addr = 6'h24;
  assign queue_bits_wb_is_ds__T_41_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_41_en = 1'h0;
  assign queue_bits_wb_is_ds__T_42_data = 1'h0;
  assign queue_bits_wb_is_ds__T_42_addr = 6'h25;
  assign queue_bits_wb_is_ds__T_42_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_42_en = 1'h0;
  assign queue_bits_wb_is_ds__T_43_data = 1'h0;
  assign queue_bits_wb_is_ds__T_43_addr = 6'h26;
  assign queue_bits_wb_is_ds__T_43_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_43_en = 1'h0;
  assign queue_bits_wb_is_ds__T_44_data = 1'h0;
  assign queue_bits_wb_is_ds__T_44_addr = 6'h27;
  assign queue_bits_wb_is_ds__T_44_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_44_en = 1'h0;
  assign queue_bits_wb_is_ds__T_45_data = 1'h0;
  assign queue_bits_wb_is_ds__T_45_addr = 6'h28;
  assign queue_bits_wb_is_ds__T_45_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_45_en = 1'h0;
  assign queue_bits_wb_is_ds__T_46_data = 1'h0;
  assign queue_bits_wb_is_ds__T_46_addr = 6'h29;
  assign queue_bits_wb_is_ds__T_46_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_46_en = 1'h0;
  assign queue_bits_wb_is_ds__T_47_data = 1'h0;
  assign queue_bits_wb_is_ds__T_47_addr = 6'h2a;
  assign queue_bits_wb_is_ds__T_47_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_47_en = 1'h0;
  assign queue_bits_wb_is_ds__T_48_data = 1'h0;
  assign queue_bits_wb_is_ds__T_48_addr = 6'h2b;
  assign queue_bits_wb_is_ds__T_48_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_48_en = 1'h0;
  assign queue_bits_wb_is_ds__T_49_data = 1'h0;
  assign queue_bits_wb_is_ds__T_49_addr = 6'h2c;
  assign queue_bits_wb_is_ds__T_49_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_49_en = 1'h0;
  assign queue_bits_wb_is_ds__T_50_data = 1'h0;
  assign queue_bits_wb_is_ds__T_50_addr = 6'h2d;
  assign queue_bits_wb_is_ds__T_50_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_50_en = 1'h0;
  assign queue_bits_wb_is_ds__T_51_data = 1'h0;
  assign queue_bits_wb_is_ds__T_51_addr = 6'h2e;
  assign queue_bits_wb_is_ds__T_51_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_51_en = 1'h0;
  assign queue_bits_wb_is_ds__T_52_data = 1'h0;
  assign queue_bits_wb_is_ds__T_52_addr = 6'h2f;
  assign queue_bits_wb_is_ds__T_52_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_52_en = 1'h0;
  assign queue_bits_wb_is_ds__T_53_data = 1'h0;
  assign queue_bits_wb_is_ds__T_53_addr = 6'h30;
  assign queue_bits_wb_is_ds__T_53_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_53_en = 1'h0;
  assign queue_bits_wb_is_ds__T_54_data = 1'h0;
  assign queue_bits_wb_is_ds__T_54_addr = 6'h31;
  assign queue_bits_wb_is_ds__T_54_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_54_en = 1'h0;
  assign queue_bits_wb_is_ds__T_55_data = 1'h0;
  assign queue_bits_wb_is_ds__T_55_addr = 6'h32;
  assign queue_bits_wb_is_ds__T_55_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_55_en = 1'h0;
  assign queue_bits_wb_is_ds__T_56_data = 1'h0;
  assign queue_bits_wb_is_ds__T_56_addr = 6'h33;
  assign queue_bits_wb_is_ds__T_56_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_56_en = 1'h0;
  assign queue_bits_wb_is_ds__T_57_data = 1'h0;
  assign queue_bits_wb_is_ds__T_57_addr = 6'h34;
  assign queue_bits_wb_is_ds__T_57_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_57_en = 1'h0;
  assign queue_bits_wb_is_ds__T_58_data = 1'h0;
  assign queue_bits_wb_is_ds__T_58_addr = 6'h35;
  assign queue_bits_wb_is_ds__T_58_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_58_en = 1'h0;
  assign queue_bits_wb_is_ds__T_59_data = 1'h0;
  assign queue_bits_wb_is_ds__T_59_addr = 6'h36;
  assign queue_bits_wb_is_ds__T_59_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_59_en = 1'h0;
  assign queue_bits_wb_is_ds__T_60_data = 1'h0;
  assign queue_bits_wb_is_ds__T_60_addr = 6'h37;
  assign queue_bits_wb_is_ds__T_60_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_60_en = 1'h0;
  assign queue_bits_wb_is_ds__T_61_data = 1'h0;
  assign queue_bits_wb_is_ds__T_61_addr = 6'h38;
  assign queue_bits_wb_is_ds__T_61_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_61_en = 1'h0;
  assign queue_bits_wb_is_ds__T_62_data = 1'h0;
  assign queue_bits_wb_is_ds__T_62_addr = 6'h39;
  assign queue_bits_wb_is_ds__T_62_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_62_en = 1'h0;
  assign queue_bits_wb_is_ds__T_63_data = 1'h0;
  assign queue_bits_wb_is_ds__T_63_addr = 6'h3a;
  assign queue_bits_wb_is_ds__T_63_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_63_en = 1'h0;
  assign queue_bits_wb_is_ds__T_64_data = 1'h0;
  assign queue_bits_wb_is_ds__T_64_addr = 6'h3b;
  assign queue_bits_wb_is_ds__T_64_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_64_en = 1'h0;
  assign queue_bits_wb_is_ds__T_65_data = 1'h0;
  assign queue_bits_wb_is_ds__T_65_addr = 6'h3c;
  assign queue_bits_wb_is_ds__T_65_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_65_en = 1'h0;
  assign queue_bits_wb_is_ds__T_66_data = 1'h0;
  assign queue_bits_wb_is_ds__T_66_addr = 6'h3d;
  assign queue_bits_wb_is_ds__T_66_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_66_en = 1'h0;
  assign queue_bits_wb_is_ds__T_67_data = 1'h0;
  assign queue_bits_wb_is_ds__T_67_addr = 6'h3e;
  assign queue_bits_wb_is_ds__T_67_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_67_en = 1'h0;
  assign queue_bits_wb_is_ds__T_68_data = 1'h0;
  assign queue_bits_wb_is_ds__T_68_addr = 6'h3f;
  assign queue_bits_wb_is_ds__T_68_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_68_en = 1'h0;
  assign queue_bits_wb_is_ds__T_70_data = 1'h0;
  assign queue_bits_wb_is_ds__T_70_addr = 6'h0;
  assign queue_bits_wb_is_ds__T_70_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_70_en = reset;
  assign queue_bits_wb_is_ds__T_71_data = 1'h0;
  assign queue_bits_wb_is_ds__T_71_addr = 6'h1;
  assign queue_bits_wb_is_ds__T_71_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_71_en = reset;
  assign queue_bits_wb_is_ds__T_72_data = 1'h0;
  assign queue_bits_wb_is_ds__T_72_addr = 6'h2;
  assign queue_bits_wb_is_ds__T_72_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_72_en = reset;
  assign queue_bits_wb_is_ds__T_73_data = 1'h0;
  assign queue_bits_wb_is_ds__T_73_addr = 6'h3;
  assign queue_bits_wb_is_ds__T_73_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_73_en = reset;
  assign queue_bits_wb_is_ds__T_74_data = 1'h0;
  assign queue_bits_wb_is_ds__T_74_addr = 6'h4;
  assign queue_bits_wb_is_ds__T_74_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_74_en = reset;
  assign queue_bits_wb_is_ds__T_75_data = 1'h0;
  assign queue_bits_wb_is_ds__T_75_addr = 6'h5;
  assign queue_bits_wb_is_ds__T_75_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_75_en = reset;
  assign queue_bits_wb_is_ds__T_76_data = 1'h0;
  assign queue_bits_wb_is_ds__T_76_addr = 6'h6;
  assign queue_bits_wb_is_ds__T_76_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_76_en = reset;
  assign queue_bits_wb_is_ds__T_77_data = 1'h0;
  assign queue_bits_wb_is_ds__T_77_addr = 6'h7;
  assign queue_bits_wb_is_ds__T_77_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_77_en = reset;
  assign queue_bits_wb_is_ds__T_78_data = 1'h0;
  assign queue_bits_wb_is_ds__T_78_addr = 6'h8;
  assign queue_bits_wb_is_ds__T_78_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_78_en = reset;
  assign queue_bits_wb_is_ds__T_79_data = 1'h0;
  assign queue_bits_wb_is_ds__T_79_addr = 6'h9;
  assign queue_bits_wb_is_ds__T_79_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_79_en = reset;
  assign queue_bits_wb_is_ds__T_80_data = 1'h0;
  assign queue_bits_wb_is_ds__T_80_addr = 6'ha;
  assign queue_bits_wb_is_ds__T_80_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_80_en = reset;
  assign queue_bits_wb_is_ds__T_81_data = 1'h0;
  assign queue_bits_wb_is_ds__T_81_addr = 6'hb;
  assign queue_bits_wb_is_ds__T_81_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_81_en = reset;
  assign queue_bits_wb_is_ds__T_82_data = 1'h0;
  assign queue_bits_wb_is_ds__T_82_addr = 6'hc;
  assign queue_bits_wb_is_ds__T_82_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_82_en = reset;
  assign queue_bits_wb_is_ds__T_83_data = 1'h0;
  assign queue_bits_wb_is_ds__T_83_addr = 6'hd;
  assign queue_bits_wb_is_ds__T_83_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_83_en = reset;
  assign queue_bits_wb_is_ds__T_84_data = 1'h0;
  assign queue_bits_wb_is_ds__T_84_addr = 6'he;
  assign queue_bits_wb_is_ds__T_84_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_84_en = reset;
  assign queue_bits_wb_is_ds__T_85_data = 1'h0;
  assign queue_bits_wb_is_ds__T_85_addr = 6'hf;
  assign queue_bits_wb_is_ds__T_85_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_85_en = reset;
  assign queue_bits_wb_is_ds__T_86_data = 1'h0;
  assign queue_bits_wb_is_ds__T_86_addr = 6'h10;
  assign queue_bits_wb_is_ds__T_86_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_86_en = reset;
  assign queue_bits_wb_is_ds__T_87_data = 1'h0;
  assign queue_bits_wb_is_ds__T_87_addr = 6'h11;
  assign queue_bits_wb_is_ds__T_87_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_87_en = reset;
  assign queue_bits_wb_is_ds__T_88_data = 1'h0;
  assign queue_bits_wb_is_ds__T_88_addr = 6'h12;
  assign queue_bits_wb_is_ds__T_88_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_88_en = reset;
  assign queue_bits_wb_is_ds__T_89_data = 1'h0;
  assign queue_bits_wb_is_ds__T_89_addr = 6'h13;
  assign queue_bits_wb_is_ds__T_89_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_89_en = reset;
  assign queue_bits_wb_is_ds__T_90_data = 1'h0;
  assign queue_bits_wb_is_ds__T_90_addr = 6'h14;
  assign queue_bits_wb_is_ds__T_90_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_90_en = reset;
  assign queue_bits_wb_is_ds__T_91_data = 1'h0;
  assign queue_bits_wb_is_ds__T_91_addr = 6'h15;
  assign queue_bits_wb_is_ds__T_91_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_91_en = reset;
  assign queue_bits_wb_is_ds__T_92_data = 1'h0;
  assign queue_bits_wb_is_ds__T_92_addr = 6'h16;
  assign queue_bits_wb_is_ds__T_92_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_92_en = reset;
  assign queue_bits_wb_is_ds__T_93_data = 1'h0;
  assign queue_bits_wb_is_ds__T_93_addr = 6'h17;
  assign queue_bits_wb_is_ds__T_93_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_93_en = reset;
  assign queue_bits_wb_is_ds__T_94_data = 1'h0;
  assign queue_bits_wb_is_ds__T_94_addr = 6'h18;
  assign queue_bits_wb_is_ds__T_94_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_94_en = reset;
  assign queue_bits_wb_is_ds__T_95_data = 1'h0;
  assign queue_bits_wb_is_ds__T_95_addr = 6'h19;
  assign queue_bits_wb_is_ds__T_95_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_95_en = reset;
  assign queue_bits_wb_is_ds__T_96_data = 1'h0;
  assign queue_bits_wb_is_ds__T_96_addr = 6'h1a;
  assign queue_bits_wb_is_ds__T_96_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_96_en = reset;
  assign queue_bits_wb_is_ds__T_97_data = 1'h0;
  assign queue_bits_wb_is_ds__T_97_addr = 6'h1b;
  assign queue_bits_wb_is_ds__T_97_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_97_en = reset;
  assign queue_bits_wb_is_ds__T_98_data = 1'h0;
  assign queue_bits_wb_is_ds__T_98_addr = 6'h1c;
  assign queue_bits_wb_is_ds__T_98_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_98_en = reset;
  assign queue_bits_wb_is_ds__T_99_data = 1'h0;
  assign queue_bits_wb_is_ds__T_99_addr = 6'h1d;
  assign queue_bits_wb_is_ds__T_99_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_99_en = reset;
  assign queue_bits_wb_is_ds__T_100_data = 1'h0;
  assign queue_bits_wb_is_ds__T_100_addr = 6'h1e;
  assign queue_bits_wb_is_ds__T_100_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_100_en = reset;
  assign queue_bits_wb_is_ds__T_101_data = 1'h0;
  assign queue_bits_wb_is_ds__T_101_addr = 6'h1f;
  assign queue_bits_wb_is_ds__T_101_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_101_en = reset;
  assign queue_bits_wb_is_ds__T_102_data = 1'h0;
  assign queue_bits_wb_is_ds__T_102_addr = 6'h20;
  assign queue_bits_wb_is_ds__T_102_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_102_en = reset;
  assign queue_bits_wb_is_ds__T_103_data = 1'h0;
  assign queue_bits_wb_is_ds__T_103_addr = 6'h21;
  assign queue_bits_wb_is_ds__T_103_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_103_en = reset;
  assign queue_bits_wb_is_ds__T_104_data = 1'h0;
  assign queue_bits_wb_is_ds__T_104_addr = 6'h22;
  assign queue_bits_wb_is_ds__T_104_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_104_en = reset;
  assign queue_bits_wb_is_ds__T_105_data = 1'h0;
  assign queue_bits_wb_is_ds__T_105_addr = 6'h23;
  assign queue_bits_wb_is_ds__T_105_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_105_en = reset;
  assign queue_bits_wb_is_ds__T_106_data = 1'h0;
  assign queue_bits_wb_is_ds__T_106_addr = 6'h24;
  assign queue_bits_wb_is_ds__T_106_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_106_en = reset;
  assign queue_bits_wb_is_ds__T_107_data = 1'h0;
  assign queue_bits_wb_is_ds__T_107_addr = 6'h25;
  assign queue_bits_wb_is_ds__T_107_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_107_en = reset;
  assign queue_bits_wb_is_ds__T_108_data = 1'h0;
  assign queue_bits_wb_is_ds__T_108_addr = 6'h26;
  assign queue_bits_wb_is_ds__T_108_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_108_en = reset;
  assign queue_bits_wb_is_ds__T_109_data = 1'h0;
  assign queue_bits_wb_is_ds__T_109_addr = 6'h27;
  assign queue_bits_wb_is_ds__T_109_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_109_en = reset;
  assign queue_bits_wb_is_ds__T_110_data = 1'h0;
  assign queue_bits_wb_is_ds__T_110_addr = 6'h28;
  assign queue_bits_wb_is_ds__T_110_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_110_en = reset;
  assign queue_bits_wb_is_ds__T_111_data = 1'h0;
  assign queue_bits_wb_is_ds__T_111_addr = 6'h29;
  assign queue_bits_wb_is_ds__T_111_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_111_en = reset;
  assign queue_bits_wb_is_ds__T_112_data = 1'h0;
  assign queue_bits_wb_is_ds__T_112_addr = 6'h2a;
  assign queue_bits_wb_is_ds__T_112_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_112_en = reset;
  assign queue_bits_wb_is_ds__T_113_data = 1'h0;
  assign queue_bits_wb_is_ds__T_113_addr = 6'h2b;
  assign queue_bits_wb_is_ds__T_113_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_113_en = reset;
  assign queue_bits_wb_is_ds__T_114_data = 1'h0;
  assign queue_bits_wb_is_ds__T_114_addr = 6'h2c;
  assign queue_bits_wb_is_ds__T_114_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_114_en = reset;
  assign queue_bits_wb_is_ds__T_115_data = 1'h0;
  assign queue_bits_wb_is_ds__T_115_addr = 6'h2d;
  assign queue_bits_wb_is_ds__T_115_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_115_en = reset;
  assign queue_bits_wb_is_ds__T_116_data = 1'h0;
  assign queue_bits_wb_is_ds__T_116_addr = 6'h2e;
  assign queue_bits_wb_is_ds__T_116_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_116_en = reset;
  assign queue_bits_wb_is_ds__T_117_data = 1'h0;
  assign queue_bits_wb_is_ds__T_117_addr = 6'h2f;
  assign queue_bits_wb_is_ds__T_117_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_117_en = reset;
  assign queue_bits_wb_is_ds__T_118_data = 1'h0;
  assign queue_bits_wb_is_ds__T_118_addr = 6'h30;
  assign queue_bits_wb_is_ds__T_118_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_118_en = reset;
  assign queue_bits_wb_is_ds__T_119_data = 1'h0;
  assign queue_bits_wb_is_ds__T_119_addr = 6'h31;
  assign queue_bits_wb_is_ds__T_119_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_119_en = reset;
  assign queue_bits_wb_is_ds__T_120_data = 1'h0;
  assign queue_bits_wb_is_ds__T_120_addr = 6'h32;
  assign queue_bits_wb_is_ds__T_120_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_120_en = reset;
  assign queue_bits_wb_is_ds__T_121_data = 1'h0;
  assign queue_bits_wb_is_ds__T_121_addr = 6'h33;
  assign queue_bits_wb_is_ds__T_121_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_121_en = reset;
  assign queue_bits_wb_is_ds__T_122_data = 1'h0;
  assign queue_bits_wb_is_ds__T_122_addr = 6'h34;
  assign queue_bits_wb_is_ds__T_122_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_122_en = reset;
  assign queue_bits_wb_is_ds__T_123_data = 1'h0;
  assign queue_bits_wb_is_ds__T_123_addr = 6'h35;
  assign queue_bits_wb_is_ds__T_123_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_123_en = reset;
  assign queue_bits_wb_is_ds__T_124_data = 1'h0;
  assign queue_bits_wb_is_ds__T_124_addr = 6'h36;
  assign queue_bits_wb_is_ds__T_124_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_124_en = reset;
  assign queue_bits_wb_is_ds__T_125_data = 1'h0;
  assign queue_bits_wb_is_ds__T_125_addr = 6'h37;
  assign queue_bits_wb_is_ds__T_125_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_125_en = reset;
  assign queue_bits_wb_is_ds__T_126_data = 1'h0;
  assign queue_bits_wb_is_ds__T_126_addr = 6'h38;
  assign queue_bits_wb_is_ds__T_126_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_126_en = reset;
  assign queue_bits_wb_is_ds__T_127_data = 1'h0;
  assign queue_bits_wb_is_ds__T_127_addr = 6'h39;
  assign queue_bits_wb_is_ds__T_127_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_127_en = reset;
  assign queue_bits_wb_is_ds__T_128_data = 1'h0;
  assign queue_bits_wb_is_ds__T_128_addr = 6'h3a;
  assign queue_bits_wb_is_ds__T_128_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_128_en = reset;
  assign queue_bits_wb_is_ds__T_129_data = 1'h0;
  assign queue_bits_wb_is_ds__T_129_addr = 6'h3b;
  assign queue_bits_wb_is_ds__T_129_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_129_en = reset;
  assign queue_bits_wb_is_ds__T_130_data = 1'h0;
  assign queue_bits_wb_is_ds__T_130_addr = 6'h3c;
  assign queue_bits_wb_is_ds__T_130_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_130_en = reset;
  assign queue_bits_wb_is_ds__T_131_data = 1'h0;
  assign queue_bits_wb_is_ds__T_131_addr = 6'h3d;
  assign queue_bits_wb_is_ds__T_131_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_131_en = reset;
  assign queue_bits_wb_is_ds__T_132_data = 1'h0;
  assign queue_bits_wb_is_ds__T_132_addr = 6'h3e;
  assign queue_bits_wb_is_ds__T_132_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_132_en = reset;
  assign queue_bits_wb_is_ds__T_133_data = 1'h0;
  assign queue_bits_wb_is_ds__T_133_addr = 6'h3f;
  assign queue_bits_wb_is_ds__T_133_mask = 1'h0;
  assign queue_bits_wb_is_ds__T_133_en = reset;
  assign queue_bits_wb_is_ds_q_head_w_data = 1'h0;
  assign queue_bits_wb_is_ds_q_head_w_addr = head;
  assign queue_bits_wb_is_ds_q_head_w_mask = 1'h0;
  assign queue_bits_wb_is_ds_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_is_br_q_head_r_addr = head;
  assign queue_bits_wb_is_br_q_head_r_data = queue_bits_wb_is_br[queue_bits_wb_is_br_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_is_br__T_3_data = io_enq_0_bits_data_wb_is_br;
  assign queue_bits_wb_is_br__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_is_br__T_3_mask = 1'h1;
  assign queue_bits_wb_is_br__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_is_br__T_4_data = io_enq_1_bits_data_wb_is_br;
  assign queue_bits_wb_is_br__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_is_br__T_4_mask = 1'h1;
  assign queue_bits_wb_is_br__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_is_br__T_5_data = 1'h0;
  assign queue_bits_wb_is_br__T_5_addr = 6'h0;
  assign queue_bits_wb_is_br__T_5_mask = 1'h0;
  assign queue_bits_wb_is_br__T_5_en = 1'h0;
  assign queue_bits_wb_is_br__T_6_data = 1'h0;
  assign queue_bits_wb_is_br__T_6_addr = 6'h1;
  assign queue_bits_wb_is_br__T_6_mask = 1'h0;
  assign queue_bits_wb_is_br__T_6_en = 1'h0;
  assign queue_bits_wb_is_br__T_7_data = 1'h0;
  assign queue_bits_wb_is_br__T_7_addr = 6'h2;
  assign queue_bits_wb_is_br__T_7_mask = 1'h0;
  assign queue_bits_wb_is_br__T_7_en = 1'h0;
  assign queue_bits_wb_is_br__T_8_data = 1'h0;
  assign queue_bits_wb_is_br__T_8_addr = 6'h3;
  assign queue_bits_wb_is_br__T_8_mask = 1'h0;
  assign queue_bits_wb_is_br__T_8_en = 1'h0;
  assign queue_bits_wb_is_br__T_9_data = 1'h0;
  assign queue_bits_wb_is_br__T_9_addr = 6'h4;
  assign queue_bits_wb_is_br__T_9_mask = 1'h0;
  assign queue_bits_wb_is_br__T_9_en = 1'h0;
  assign queue_bits_wb_is_br__T_10_data = 1'h0;
  assign queue_bits_wb_is_br__T_10_addr = 6'h5;
  assign queue_bits_wb_is_br__T_10_mask = 1'h0;
  assign queue_bits_wb_is_br__T_10_en = 1'h0;
  assign queue_bits_wb_is_br__T_11_data = 1'h0;
  assign queue_bits_wb_is_br__T_11_addr = 6'h6;
  assign queue_bits_wb_is_br__T_11_mask = 1'h0;
  assign queue_bits_wb_is_br__T_11_en = 1'h0;
  assign queue_bits_wb_is_br__T_12_data = 1'h0;
  assign queue_bits_wb_is_br__T_12_addr = 6'h7;
  assign queue_bits_wb_is_br__T_12_mask = 1'h0;
  assign queue_bits_wb_is_br__T_12_en = 1'h0;
  assign queue_bits_wb_is_br__T_13_data = 1'h0;
  assign queue_bits_wb_is_br__T_13_addr = 6'h8;
  assign queue_bits_wb_is_br__T_13_mask = 1'h0;
  assign queue_bits_wb_is_br__T_13_en = 1'h0;
  assign queue_bits_wb_is_br__T_14_data = 1'h0;
  assign queue_bits_wb_is_br__T_14_addr = 6'h9;
  assign queue_bits_wb_is_br__T_14_mask = 1'h0;
  assign queue_bits_wb_is_br__T_14_en = 1'h0;
  assign queue_bits_wb_is_br__T_15_data = 1'h0;
  assign queue_bits_wb_is_br__T_15_addr = 6'ha;
  assign queue_bits_wb_is_br__T_15_mask = 1'h0;
  assign queue_bits_wb_is_br__T_15_en = 1'h0;
  assign queue_bits_wb_is_br__T_16_data = 1'h0;
  assign queue_bits_wb_is_br__T_16_addr = 6'hb;
  assign queue_bits_wb_is_br__T_16_mask = 1'h0;
  assign queue_bits_wb_is_br__T_16_en = 1'h0;
  assign queue_bits_wb_is_br__T_17_data = 1'h0;
  assign queue_bits_wb_is_br__T_17_addr = 6'hc;
  assign queue_bits_wb_is_br__T_17_mask = 1'h0;
  assign queue_bits_wb_is_br__T_17_en = 1'h0;
  assign queue_bits_wb_is_br__T_18_data = 1'h0;
  assign queue_bits_wb_is_br__T_18_addr = 6'hd;
  assign queue_bits_wb_is_br__T_18_mask = 1'h0;
  assign queue_bits_wb_is_br__T_18_en = 1'h0;
  assign queue_bits_wb_is_br__T_19_data = 1'h0;
  assign queue_bits_wb_is_br__T_19_addr = 6'he;
  assign queue_bits_wb_is_br__T_19_mask = 1'h0;
  assign queue_bits_wb_is_br__T_19_en = 1'h0;
  assign queue_bits_wb_is_br__T_20_data = 1'h0;
  assign queue_bits_wb_is_br__T_20_addr = 6'hf;
  assign queue_bits_wb_is_br__T_20_mask = 1'h0;
  assign queue_bits_wb_is_br__T_20_en = 1'h0;
  assign queue_bits_wb_is_br__T_21_data = 1'h0;
  assign queue_bits_wb_is_br__T_21_addr = 6'h10;
  assign queue_bits_wb_is_br__T_21_mask = 1'h0;
  assign queue_bits_wb_is_br__T_21_en = 1'h0;
  assign queue_bits_wb_is_br__T_22_data = 1'h0;
  assign queue_bits_wb_is_br__T_22_addr = 6'h11;
  assign queue_bits_wb_is_br__T_22_mask = 1'h0;
  assign queue_bits_wb_is_br__T_22_en = 1'h0;
  assign queue_bits_wb_is_br__T_23_data = 1'h0;
  assign queue_bits_wb_is_br__T_23_addr = 6'h12;
  assign queue_bits_wb_is_br__T_23_mask = 1'h0;
  assign queue_bits_wb_is_br__T_23_en = 1'h0;
  assign queue_bits_wb_is_br__T_24_data = 1'h0;
  assign queue_bits_wb_is_br__T_24_addr = 6'h13;
  assign queue_bits_wb_is_br__T_24_mask = 1'h0;
  assign queue_bits_wb_is_br__T_24_en = 1'h0;
  assign queue_bits_wb_is_br__T_25_data = 1'h0;
  assign queue_bits_wb_is_br__T_25_addr = 6'h14;
  assign queue_bits_wb_is_br__T_25_mask = 1'h0;
  assign queue_bits_wb_is_br__T_25_en = 1'h0;
  assign queue_bits_wb_is_br__T_26_data = 1'h0;
  assign queue_bits_wb_is_br__T_26_addr = 6'h15;
  assign queue_bits_wb_is_br__T_26_mask = 1'h0;
  assign queue_bits_wb_is_br__T_26_en = 1'h0;
  assign queue_bits_wb_is_br__T_27_data = 1'h0;
  assign queue_bits_wb_is_br__T_27_addr = 6'h16;
  assign queue_bits_wb_is_br__T_27_mask = 1'h0;
  assign queue_bits_wb_is_br__T_27_en = 1'h0;
  assign queue_bits_wb_is_br__T_28_data = 1'h0;
  assign queue_bits_wb_is_br__T_28_addr = 6'h17;
  assign queue_bits_wb_is_br__T_28_mask = 1'h0;
  assign queue_bits_wb_is_br__T_28_en = 1'h0;
  assign queue_bits_wb_is_br__T_29_data = 1'h0;
  assign queue_bits_wb_is_br__T_29_addr = 6'h18;
  assign queue_bits_wb_is_br__T_29_mask = 1'h0;
  assign queue_bits_wb_is_br__T_29_en = 1'h0;
  assign queue_bits_wb_is_br__T_30_data = 1'h0;
  assign queue_bits_wb_is_br__T_30_addr = 6'h19;
  assign queue_bits_wb_is_br__T_30_mask = 1'h0;
  assign queue_bits_wb_is_br__T_30_en = 1'h0;
  assign queue_bits_wb_is_br__T_31_data = 1'h0;
  assign queue_bits_wb_is_br__T_31_addr = 6'h1a;
  assign queue_bits_wb_is_br__T_31_mask = 1'h0;
  assign queue_bits_wb_is_br__T_31_en = 1'h0;
  assign queue_bits_wb_is_br__T_32_data = 1'h0;
  assign queue_bits_wb_is_br__T_32_addr = 6'h1b;
  assign queue_bits_wb_is_br__T_32_mask = 1'h0;
  assign queue_bits_wb_is_br__T_32_en = 1'h0;
  assign queue_bits_wb_is_br__T_33_data = 1'h0;
  assign queue_bits_wb_is_br__T_33_addr = 6'h1c;
  assign queue_bits_wb_is_br__T_33_mask = 1'h0;
  assign queue_bits_wb_is_br__T_33_en = 1'h0;
  assign queue_bits_wb_is_br__T_34_data = 1'h0;
  assign queue_bits_wb_is_br__T_34_addr = 6'h1d;
  assign queue_bits_wb_is_br__T_34_mask = 1'h0;
  assign queue_bits_wb_is_br__T_34_en = 1'h0;
  assign queue_bits_wb_is_br__T_35_data = 1'h0;
  assign queue_bits_wb_is_br__T_35_addr = 6'h1e;
  assign queue_bits_wb_is_br__T_35_mask = 1'h0;
  assign queue_bits_wb_is_br__T_35_en = 1'h0;
  assign queue_bits_wb_is_br__T_36_data = 1'h0;
  assign queue_bits_wb_is_br__T_36_addr = 6'h1f;
  assign queue_bits_wb_is_br__T_36_mask = 1'h0;
  assign queue_bits_wb_is_br__T_36_en = 1'h0;
  assign queue_bits_wb_is_br__T_37_data = 1'h0;
  assign queue_bits_wb_is_br__T_37_addr = 6'h20;
  assign queue_bits_wb_is_br__T_37_mask = 1'h0;
  assign queue_bits_wb_is_br__T_37_en = 1'h0;
  assign queue_bits_wb_is_br__T_38_data = 1'h0;
  assign queue_bits_wb_is_br__T_38_addr = 6'h21;
  assign queue_bits_wb_is_br__T_38_mask = 1'h0;
  assign queue_bits_wb_is_br__T_38_en = 1'h0;
  assign queue_bits_wb_is_br__T_39_data = 1'h0;
  assign queue_bits_wb_is_br__T_39_addr = 6'h22;
  assign queue_bits_wb_is_br__T_39_mask = 1'h0;
  assign queue_bits_wb_is_br__T_39_en = 1'h0;
  assign queue_bits_wb_is_br__T_40_data = 1'h0;
  assign queue_bits_wb_is_br__T_40_addr = 6'h23;
  assign queue_bits_wb_is_br__T_40_mask = 1'h0;
  assign queue_bits_wb_is_br__T_40_en = 1'h0;
  assign queue_bits_wb_is_br__T_41_data = 1'h0;
  assign queue_bits_wb_is_br__T_41_addr = 6'h24;
  assign queue_bits_wb_is_br__T_41_mask = 1'h0;
  assign queue_bits_wb_is_br__T_41_en = 1'h0;
  assign queue_bits_wb_is_br__T_42_data = 1'h0;
  assign queue_bits_wb_is_br__T_42_addr = 6'h25;
  assign queue_bits_wb_is_br__T_42_mask = 1'h0;
  assign queue_bits_wb_is_br__T_42_en = 1'h0;
  assign queue_bits_wb_is_br__T_43_data = 1'h0;
  assign queue_bits_wb_is_br__T_43_addr = 6'h26;
  assign queue_bits_wb_is_br__T_43_mask = 1'h0;
  assign queue_bits_wb_is_br__T_43_en = 1'h0;
  assign queue_bits_wb_is_br__T_44_data = 1'h0;
  assign queue_bits_wb_is_br__T_44_addr = 6'h27;
  assign queue_bits_wb_is_br__T_44_mask = 1'h0;
  assign queue_bits_wb_is_br__T_44_en = 1'h0;
  assign queue_bits_wb_is_br__T_45_data = 1'h0;
  assign queue_bits_wb_is_br__T_45_addr = 6'h28;
  assign queue_bits_wb_is_br__T_45_mask = 1'h0;
  assign queue_bits_wb_is_br__T_45_en = 1'h0;
  assign queue_bits_wb_is_br__T_46_data = 1'h0;
  assign queue_bits_wb_is_br__T_46_addr = 6'h29;
  assign queue_bits_wb_is_br__T_46_mask = 1'h0;
  assign queue_bits_wb_is_br__T_46_en = 1'h0;
  assign queue_bits_wb_is_br__T_47_data = 1'h0;
  assign queue_bits_wb_is_br__T_47_addr = 6'h2a;
  assign queue_bits_wb_is_br__T_47_mask = 1'h0;
  assign queue_bits_wb_is_br__T_47_en = 1'h0;
  assign queue_bits_wb_is_br__T_48_data = 1'h0;
  assign queue_bits_wb_is_br__T_48_addr = 6'h2b;
  assign queue_bits_wb_is_br__T_48_mask = 1'h0;
  assign queue_bits_wb_is_br__T_48_en = 1'h0;
  assign queue_bits_wb_is_br__T_49_data = 1'h0;
  assign queue_bits_wb_is_br__T_49_addr = 6'h2c;
  assign queue_bits_wb_is_br__T_49_mask = 1'h0;
  assign queue_bits_wb_is_br__T_49_en = 1'h0;
  assign queue_bits_wb_is_br__T_50_data = 1'h0;
  assign queue_bits_wb_is_br__T_50_addr = 6'h2d;
  assign queue_bits_wb_is_br__T_50_mask = 1'h0;
  assign queue_bits_wb_is_br__T_50_en = 1'h0;
  assign queue_bits_wb_is_br__T_51_data = 1'h0;
  assign queue_bits_wb_is_br__T_51_addr = 6'h2e;
  assign queue_bits_wb_is_br__T_51_mask = 1'h0;
  assign queue_bits_wb_is_br__T_51_en = 1'h0;
  assign queue_bits_wb_is_br__T_52_data = 1'h0;
  assign queue_bits_wb_is_br__T_52_addr = 6'h2f;
  assign queue_bits_wb_is_br__T_52_mask = 1'h0;
  assign queue_bits_wb_is_br__T_52_en = 1'h0;
  assign queue_bits_wb_is_br__T_53_data = 1'h0;
  assign queue_bits_wb_is_br__T_53_addr = 6'h30;
  assign queue_bits_wb_is_br__T_53_mask = 1'h0;
  assign queue_bits_wb_is_br__T_53_en = 1'h0;
  assign queue_bits_wb_is_br__T_54_data = 1'h0;
  assign queue_bits_wb_is_br__T_54_addr = 6'h31;
  assign queue_bits_wb_is_br__T_54_mask = 1'h0;
  assign queue_bits_wb_is_br__T_54_en = 1'h0;
  assign queue_bits_wb_is_br__T_55_data = 1'h0;
  assign queue_bits_wb_is_br__T_55_addr = 6'h32;
  assign queue_bits_wb_is_br__T_55_mask = 1'h0;
  assign queue_bits_wb_is_br__T_55_en = 1'h0;
  assign queue_bits_wb_is_br__T_56_data = 1'h0;
  assign queue_bits_wb_is_br__T_56_addr = 6'h33;
  assign queue_bits_wb_is_br__T_56_mask = 1'h0;
  assign queue_bits_wb_is_br__T_56_en = 1'h0;
  assign queue_bits_wb_is_br__T_57_data = 1'h0;
  assign queue_bits_wb_is_br__T_57_addr = 6'h34;
  assign queue_bits_wb_is_br__T_57_mask = 1'h0;
  assign queue_bits_wb_is_br__T_57_en = 1'h0;
  assign queue_bits_wb_is_br__T_58_data = 1'h0;
  assign queue_bits_wb_is_br__T_58_addr = 6'h35;
  assign queue_bits_wb_is_br__T_58_mask = 1'h0;
  assign queue_bits_wb_is_br__T_58_en = 1'h0;
  assign queue_bits_wb_is_br__T_59_data = 1'h0;
  assign queue_bits_wb_is_br__T_59_addr = 6'h36;
  assign queue_bits_wb_is_br__T_59_mask = 1'h0;
  assign queue_bits_wb_is_br__T_59_en = 1'h0;
  assign queue_bits_wb_is_br__T_60_data = 1'h0;
  assign queue_bits_wb_is_br__T_60_addr = 6'h37;
  assign queue_bits_wb_is_br__T_60_mask = 1'h0;
  assign queue_bits_wb_is_br__T_60_en = 1'h0;
  assign queue_bits_wb_is_br__T_61_data = 1'h0;
  assign queue_bits_wb_is_br__T_61_addr = 6'h38;
  assign queue_bits_wb_is_br__T_61_mask = 1'h0;
  assign queue_bits_wb_is_br__T_61_en = 1'h0;
  assign queue_bits_wb_is_br__T_62_data = 1'h0;
  assign queue_bits_wb_is_br__T_62_addr = 6'h39;
  assign queue_bits_wb_is_br__T_62_mask = 1'h0;
  assign queue_bits_wb_is_br__T_62_en = 1'h0;
  assign queue_bits_wb_is_br__T_63_data = 1'h0;
  assign queue_bits_wb_is_br__T_63_addr = 6'h3a;
  assign queue_bits_wb_is_br__T_63_mask = 1'h0;
  assign queue_bits_wb_is_br__T_63_en = 1'h0;
  assign queue_bits_wb_is_br__T_64_data = 1'h0;
  assign queue_bits_wb_is_br__T_64_addr = 6'h3b;
  assign queue_bits_wb_is_br__T_64_mask = 1'h0;
  assign queue_bits_wb_is_br__T_64_en = 1'h0;
  assign queue_bits_wb_is_br__T_65_data = 1'h0;
  assign queue_bits_wb_is_br__T_65_addr = 6'h3c;
  assign queue_bits_wb_is_br__T_65_mask = 1'h0;
  assign queue_bits_wb_is_br__T_65_en = 1'h0;
  assign queue_bits_wb_is_br__T_66_data = 1'h0;
  assign queue_bits_wb_is_br__T_66_addr = 6'h3d;
  assign queue_bits_wb_is_br__T_66_mask = 1'h0;
  assign queue_bits_wb_is_br__T_66_en = 1'h0;
  assign queue_bits_wb_is_br__T_67_data = 1'h0;
  assign queue_bits_wb_is_br__T_67_addr = 6'h3e;
  assign queue_bits_wb_is_br__T_67_mask = 1'h0;
  assign queue_bits_wb_is_br__T_67_en = 1'h0;
  assign queue_bits_wb_is_br__T_68_data = 1'h0;
  assign queue_bits_wb_is_br__T_68_addr = 6'h3f;
  assign queue_bits_wb_is_br__T_68_mask = 1'h0;
  assign queue_bits_wb_is_br__T_68_en = 1'h0;
  assign queue_bits_wb_is_br__T_70_data = 1'h0;
  assign queue_bits_wb_is_br__T_70_addr = 6'h0;
  assign queue_bits_wb_is_br__T_70_mask = 1'h0;
  assign queue_bits_wb_is_br__T_70_en = reset;
  assign queue_bits_wb_is_br__T_71_data = 1'h0;
  assign queue_bits_wb_is_br__T_71_addr = 6'h1;
  assign queue_bits_wb_is_br__T_71_mask = 1'h0;
  assign queue_bits_wb_is_br__T_71_en = reset;
  assign queue_bits_wb_is_br__T_72_data = 1'h0;
  assign queue_bits_wb_is_br__T_72_addr = 6'h2;
  assign queue_bits_wb_is_br__T_72_mask = 1'h0;
  assign queue_bits_wb_is_br__T_72_en = reset;
  assign queue_bits_wb_is_br__T_73_data = 1'h0;
  assign queue_bits_wb_is_br__T_73_addr = 6'h3;
  assign queue_bits_wb_is_br__T_73_mask = 1'h0;
  assign queue_bits_wb_is_br__T_73_en = reset;
  assign queue_bits_wb_is_br__T_74_data = 1'h0;
  assign queue_bits_wb_is_br__T_74_addr = 6'h4;
  assign queue_bits_wb_is_br__T_74_mask = 1'h0;
  assign queue_bits_wb_is_br__T_74_en = reset;
  assign queue_bits_wb_is_br__T_75_data = 1'h0;
  assign queue_bits_wb_is_br__T_75_addr = 6'h5;
  assign queue_bits_wb_is_br__T_75_mask = 1'h0;
  assign queue_bits_wb_is_br__T_75_en = reset;
  assign queue_bits_wb_is_br__T_76_data = 1'h0;
  assign queue_bits_wb_is_br__T_76_addr = 6'h6;
  assign queue_bits_wb_is_br__T_76_mask = 1'h0;
  assign queue_bits_wb_is_br__T_76_en = reset;
  assign queue_bits_wb_is_br__T_77_data = 1'h0;
  assign queue_bits_wb_is_br__T_77_addr = 6'h7;
  assign queue_bits_wb_is_br__T_77_mask = 1'h0;
  assign queue_bits_wb_is_br__T_77_en = reset;
  assign queue_bits_wb_is_br__T_78_data = 1'h0;
  assign queue_bits_wb_is_br__T_78_addr = 6'h8;
  assign queue_bits_wb_is_br__T_78_mask = 1'h0;
  assign queue_bits_wb_is_br__T_78_en = reset;
  assign queue_bits_wb_is_br__T_79_data = 1'h0;
  assign queue_bits_wb_is_br__T_79_addr = 6'h9;
  assign queue_bits_wb_is_br__T_79_mask = 1'h0;
  assign queue_bits_wb_is_br__T_79_en = reset;
  assign queue_bits_wb_is_br__T_80_data = 1'h0;
  assign queue_bits_wb_is_br__T_80_addr = 6'ha;
  assign queue_bits_wb_is_br__T_80_mask = 1'h0;
  assign queue_bits_wb_is_br__T_80_en = reset;
  assign queue_bits_wb_is_br__T_81_data = 1'h0;
  assign queue_bits_wb_is_br__T_81_addr = 6'hb;
  assign queue_bits_wb_is_br__T_81_mask = 1'h0;
  assign queue_bits_wb_is_br__T_81_en = reset;
  assign queue_bits_wb_is_br__T_82_data = 1'h0;
  assign queue_bits_wb_is_br__T_82_addr = 6'hc;
  assign queue_bits_wb_is_br__T_82_mask = 1'h0;
  assign queue_bits_wb_is_br__T_82_en = reset;
  assign queue_bits_wb_is_br__T_83_data = 1'h0;
  assign queue_bits_wb_is_br__T_83_addr = 6'hd;
  assign queue_bits_wb_is_br__T_83_mask = 1'h0;
  assign queue_bits_wb_is_br__T_83_en = reset;
  assign queue_bits_wb_is_br__T_84_data = 1'h0;
  assign queue_bits_wb_is_br__T_84_addr = 6'he;
  assign queue_bits_wb_is_br__T_84_mask = 1'h0;
  assign queue_bits_wb_is_br__T_84_en = reset;
  assign queue_bits_wb_is_br__T_85_data = 1'h0;
  assign queue_bits_wb_is_br__T_85_addr = 6'hf;
  assign queue_bits_wb_is_br__T_85_mask = 1'h0;
  assign queue_bits_wb_is_br__T_85_en = reset;
  assign queue_bits_wb_is_br__T_86_data = 1'h0;
  assign queue_bits_wb_is_br__T_86_addr = 6'h10;
  assign queue_bits_wb_is_br__T_86_mask = 1'h0;
  assign queue_bits_wb_is_br__T_86_en = reset;
  assign queue_bits_wb_is_br__T_87_data = 1'h0;
  assign queue_bits_wb_is_br__T_87_addr = 6'h11;
  assign queue_bits_wb_is_br__T_87_mask = 1'h0;
  assign queue_bits_wb_is_br__T_87_en = reset;
  assign queue_bits_wb_is_br__T_88_data = 1'h0;
  assign queue_bits_wb_is_br__T_88_addr = 6'h12;
  assign queue_bits_wb_is_br__T_88_mask = 1'h0;
  assign queue_bits_wb_is_br__T_88_en = reset;
  assign queue_bits_wb_is_br__T_89_data = 1'h0;
  assign queue_bits_wb_is_br__T_89_addr = 6'h13;
  assign queue_bits_wb_is_br__T_89_mask = 1'h0;
  assign queue_bits_wb_is_br__T_89_en = reset;
  assign queue_bits_wb_is_br__T_90_data = 1'h0;
  assign queue_bits_wb_is_br__T_90_addr = 6'h14;
  assign queue_bits_wb_is_br__T_90_mask = 1'h0;
  assign queue_bits_wb_is_br__T_90_en = reset;
  assign queue_bits_wb_is_br__T_91_data = 1'h0;
  assign queue_bits_wb_is_br__T_91_addr = 6'h15;
  assign queue_bits_wb_is_br__T_91_mask = 1'h0;
  assign queue_bits_wb_is_br__T_91_en = reset;
  assign queue_bits_wb_is_br__T_92_data = 1'h0;
  assign queue_bits_wb_is_br__T_92_addr = 6'h16;
  assign queue_bits_wb_is_br__T_92_mask = 1'h0;
  assign queue_bits_wb_is_br__T_92_en = reset;
  assign queue_bits_wb_is_br__T_93_data = 1'h0;
  assign queue_bits_wb_is_br__T_93_addr = 6'h17;
  assign queue_bits_wb_is_br__T_93_mask = 1'h0;
  assign queue_bits_wb_is_br__T_93_en = reset;
  assign queue_bits_wb_is_br__T_94_data = 1'h0;
  assign queue_bits_wb_is_br__T_94_addr = 6'h18;
  assign queue_bits_wb_is_br__T_94_mask = 1'h0;
  assign queue_bits_wb_is_br__T_94_en = reset;
  assign queue_bits_wb_is_br__T_95_data = 1'h0;
  assign queue_bits_wb_is_br__T_95_addr = 6'h19;
  assign queue_bits_wb_is_br__T_95_mask = 1'h0;
  assign queue_bits_wb_is_br__T_95_en = reset;
  assign queue_bits_wb_is_br__T_96_data = 1'h0;
  assign queue_bits_wb_is_br__T_96_addr = 6'h1a;
  assign queue_bits_wb_is_br__T_96_mask = 1'h0;
  assign queue_bits_wb_is_br__T_96_en = reset;
  assign queue_bits_wb_is_br__T_97_data = 1'h0;
  assign queue_bits_wb_is_br__T_97_addr = 6'h1b;
  assign queue_bits_wb_is_br__T_97_mask = 1'h0;
  assign queue_bits_wb_is_br__T_97_en = reset;
  assign queue_bits_wb_is_br__T_98_data = 1'h0;
  assign queue_bits_wb_is_br__T_98_addr = 6'h1c;
  assign queue_bits_wb_is_br__T_98_mask = 1'h0;
  assign queue_bits_wb_is_br__T_98_en = reset;
  assign queue_bits_wb_is_br__T_99_data = 1'h0;
  assign queue_bits_wb_is_br__T_99_addr = 6'h1d;
  assign queue_bits_wb_is_br__T_99_mask = 1'h0;
  assign queue_bits_wb_is_br__T_99_en = reset;
  assign queue_bits_wb_is_br__T_100_data = 1'h0;
  assign queue_bits_wb_is_br__T_100_addr = 6'h1e;
  assign queue_bits_wb_is_br__T_100_mask = 1'h0;
  assign queue_bits_wb_is_br__T_100_en = reset;
  assign queue_bits_wb_is_br__T_101_data = 1'h0;
  assign queue_bits_wb_is_br__T_101_addr = 6'h1f;
  assign queue_bits_wb_is_br__T_101_mask = 1'h0;
  assign queue_bits_wb_is_br__T_101_en = reset;
  assign queue_bits_wb_is_br__T_102_data = 1'h0;
  assign queue_bits_wb_is_br__T_102_addr = 6'h20;
  assign queue_bits_wb_is_br__T_102_mask = 1'h0;
  assign queue_bits_wb_is_br__T_102_en = reset;
  assign queue_bits_wb_is_br__T_103_data = 1'h0;
  assign queue_bits_wb_is_br__T_103_addr = 6'h21;
  assign queue_bits_wb_is_br__T_103_mask = 1'h0;
  assign queue_bits_wb_is_br__T_103_en = reset;
  assign queue_bits_wb_is_br__T_104_data = 1'h0;
  assign queue_bits_wb_is_br__T_104_addr = 6'h22;
  assign queue_bits_wb_is_br__T_104_mask = 1'h0;
  assign queue_bits_wb_is_br__T_104_en = reset;
  assign queue_bits_wb_is_br__T_105_data = 1'h0;
  assign queue_bits_wb_is_br__T_105_addr = 6'h23;
  assign queue_bits_wb_is_br__T_105_mask = 1'h0;
  assign queue_bits_wb_is_br__T_105_en = reset;
  assign queue_bits_wb_is_br__T_106_data = 1'h0;
  assign queue_bits_wb_is_br__T_106_addr = 6'h24;
  assign queue_bits_wb_is_br__T_106_mask = 1'h0;
  assign queue_bits_wb_is_br__T_106_en = reset;
  assign queue_bits_wb_is_br__T_107_data = 1'h0;
  assign queue_bits_wb_is_br__T_107_addr = 6'h25;
  assign queue_bits_wb_is_br__T_107_mask = 1'h0;
  assign queue_bits_wb_is_br__T_107_en = reset;
  assign queue_bits_wb_is_br__T_108_data = 1'h0;
  assign queue_bits_wb_is_br__T_108_addr = 6'h26;
  assign queue_bits_wb_is_br__T_108_mask = 1'h0;
  assign queue_bits_wb_is_br__T_108_en = reset;
  assign queue_bits_wb_is_br__T_109_data = 1'h0;
  assign queue_bits_wb_is_br__T_109_addr = 6'h27;
  assign queue_bits_wb_is_br__T_109_mask = 1'h0;
  assign queue_bits_wb_is_br__T_109_en = reset;
  assign queue_bits_wb_is_br__T_110_data = 1'h0;
  assign queue_bits_wb_is_br__T_110_addr = 6'h28;
  assign queue_bits_wb_is_br__T_110_mask = 1'h0;
  assign queue_bits_wb_is_br__T_110_en = reset;
  assign queue_bits_wb_is_br__T_111_data = 1'h0;
  assign queue_bits_wb_is_br__T_111_addr = 6'h29;
  assign queue_bits_wb_is_br__T_111_mask = 1'h0;
  assign queue_bits_wb_is_br__T_111_en = reset;
  assign queue_bits_wb_is_br__T_112_data = 1'h0;
  assign queue_bits_wb_is_br__T_112_addr = 6'h2a;
  assign queue_bits_wb_is_br__T_112_mask = 1'h0;
  assign queue_bits_wb_is_br__T_112_en = reset;
  assign queue_bits_wb_is_br__T_113_data = 1'h0;
  assign queue_bits_wb_is_br__T_113_addr = 6'h2b;
  assign queue_bits_wb_is_br__T_113_mask = 1'h0;
  assign queue_bits_wb_is_br__T_113_en = reset;
  assign queue_bits_wb_is_br__T_114_data = 1'h0;
  assign queue_bits_wb_is_br__T_114_addr = 6'h2c;
  assign queue_bits_wb_is_br__T_114_mask = 1'h0;
  assign queue_bits_wb_is_br__T_114_en = reset;
  assign queue_bits_wb_is_br__T_115_data = 1'h0;
  assign queue_bits_wb_is_br__T_115_addr = 6'h2d;
  assign queue_bits_wb_is_br__T_115_mask = 1'h0;
  assign queue_bits_wb_is_br__T_115_en = reset;
  assign queue_bits_wb_is_br__T_116_data = 1'h0;
  assign queue_bits_wb_is_br__T_116_addr = 6'h2e;
  assign queue_bits_wb_is_br__T_116_mask = 1'h0;
  assign queue_bits_wb_is_br__T_116_en = reset;
  assign queue_bits_wb_is_br__T_117_data = 1'h0;
  assign queue_bits_wb_is_br__T_117_addr = 6'h2f;
  assign queue_bits_wb_is_br__T_117_mask = 1'h0;
  assign queue_bits_wb_is_br__T_117_en = reset;
  assign queue_bits_wb_is_br__T_118_data = 1'h0;
  assign queue_bits_wb_is_br__T_118_addr = 6'h30;
  assign queue_bits_wb_is_br__T_118_mask = 1'h0;
  assign queue_bits_wb_is_br__T_118_en = reset;
  assign queue_bits_wb_is_br__T_119_data = 1'h0;
  assign queue_bits_wb_is_br__T_119_addr = 6'h31;
  assign queue_bits_wb_is_br__T_119_mask = 1'h0;
  assign queue_bits_wb_is_br__T_119_en = reset;
  assign queue_bits_wb_is_br__T_120_data = 1'h0;
  assign queue_bits_wb_is_br__T_120_addr = 6'h32;
  assign queue_bits_wb_is_br__T_120_mask = 1'h0;
  assign queue_bits_wb_is_br__T_120_en = reset;
  assign queue_bits_wb_is_br__T_121_data = 1'h0;
  assign queue_bits_wb_is_br__T_121_addr = 6'h33;
  assign queue_bits_wb_is_br__T_121_mask = 1'h0;
  assign queue_bits_wb_is_br__T_121_en = reset;
  assign queue_bits_wb_is_br__T_122_data = 1'h0;
  assign queue_bits_wb_is_br__T_122_addr = 6'h34;
  assign queue_bits_wb_is_br__T_122_mask = 1'h0;
  assign queue_bits_wb_is_br__T_122_en = reset;
  assign queue_bits_wb_is_br__T_123_data = 1'h0;
  assign queue_bits_wb_is_br__T_123_addr = 6'h35;
  assign queue_bits_wb_is_br__T_123_mask = 1'h0;
  assign queue_bits_wb_is_br__T_123_en = reset;
  assign queue_bits_wb_is_br__T_124_data = 1'h0;
  assign queue_bits_wb_is_br__T_124_addr = 6'h36;
  assign queue_bits_wb_is_br__T_124_mask = 1'h0;
  assign queue_bits_wb_is_br__T_124_en = reset;
  assign queue_bits_wb_is_br__T_125_data = 1'h0;
  assign queue_bits_wb_is_br__T_125_addr = 6'h37;
  assign queue_bits_wb_is_br__T_125_mask = 1'h0;
  assign queue_bits_wb_is_br__T_125_en = reset;
  assign queue_bits_wb_is_br__T_126_data = 1'h0;
  assign queue_bits_wb_is_br__T_126_addr = 6'h38;
  assign queue_bits_wb_is_br__T_126_mask = 1'h0;
  assign queue_bits_wb_is_br__T_126_en = reset;
  assign queue_bits_wb_is_br__T_127_data = 1'h0;
  assign queue_bits_wb_is_br__T_127_addr = 6'h39;
  assign queue_bits_wb_is_br__T_127_mask = 1'h0;
  assign queue_bits_wb_is_br__T_127_en = reset;
  assign queue_bits_wb_is_br__T_128_data = 1'h0;
  assign queue_bits_wb_is_br__T_128_addr = 6'h3a;
  assign queue_bits_wb_is_br__T_128_mask = 1'h0;
  assign queue_bits_wb_is_br__T_128_en = reset;
  assign queue_bits_wb_is_br__T_129_data = 1'h0;
  assign queue_bits_wb_is_br__T_129_addr = 6'h3b;
  assign queue_bits_wb_is_br__T_129_mask = 1'h0;
  assign queue_bits_wb_is_br__T_129_en = reset;
  assign queue_bits_wb_is_br__T_130_data = 1'h0;
  assign queue_bits_wb_is_br__T_130_addr = 6'h3c;
  assign queue_bits_wb_is_br__T_130_mask = 1'h0;
  assign queue_bits_wb_is_br__T_130_en = reset;
  assign queue_bits_wb_is_br__T_131_data = 1'h0;
  assign queue_bits_wb_is_br__T_131_addr = 6'h3d;
  assign queue_bits_wb_is_br__T_131_mask = 1'h0;
  assign queue_bits_wb_is_br__T_131_en = reset;
  assign queue_bits_wb_is_br__T_132_data = 1'h0;
  assign queue_bits_wb_is_br__T_132_addr = 6'h3e;
  assign queue_bits_wb_is_br__T_132_mask = 1'h0;
  assign queue_bits_wb_is_br__T_132_en = reset;
  assign queue_bits_wb_is_br__T_133_data = 1'h0;
  assign queue_bits_wb_is_br__T_133_addr = 6'h3f;
  assign queue_bits_wb_is_br__T_133_mask = 1'h0;
  assign queue_bits_wb_is_br__T_133_en = reset;
  assign queue_bits_wb_is_br_q_head_w_data = 1'h0;
  assign queue_bits_wb_is_br_q_head_w_addr = head;
  assign queue_bits_wb_is_br_q_head_w_mask = 1'h0;
  assign queue_bits_wb_is_br_q_head_w_en = io_deq_valid;
  assign queue_bits_wb_npc_q_head_r_addr = head;
  assign queue_bits_wb_npc_q_head_r_data = queue_bits_wb_npc[queue_bits_wb_npc_q_head_r_addr]; // @[utils.scala 30:18]
  assign queue_bits_wb_npc__T_3_data = io_enq_0_bits_data_wb_npc;
  assign queue_bits_wb_npc__T_3_addr = io_enq_0_bits_id;
  assign queue_bits_wb_npc__T_3_mask = 1'h1;
  assign queue_bits_wb_npc__T_3_en = io_enq_0_valid;
  assign queue_bits_wb_npc__T_4_data = io_enq_1_bits_data_wb_npc;
  assign queue_bits_wb_npc__T_4_addr = io_enq_1_bits_id;
  assign queue_bits_wb_npc__T_4_mask = 1'h1;
  assign queue_bits_wb_npc__T_4_en = io_enq_1_valid;
  assign queue_bits_wb_npc__T_5_data = 32'h0;
  assign queue_bits_wb_npc__T_5_addr = 6'h0;
  assign queue_bits_wb_npc__T_5_mask = 1'h0;
  assign queue_bits_wb_npc__T_5_en = 1'h0;
  assign queue_bits_wb_npc__T_6_data = 32'h0;
  assign queue_bits_wb_npc__T_6_addr = 6'h1;
  assign queue_bits_wb_npc__T_6_mask = 1'h0;
  assign queue_bits_wb_npc__T_6_en = 1'h0;
  assign queue_bits_wb_npc__T_7_data = 32'h0;
  assign queue_bits_wb_npc__T_7_addr = 6'h2;
  assign queue_bits_wb_npc__T_7_mask = 1'h0;
  assign queue_bits_wb_npc__T_7_en = 1'h0;
  assign queue_bits_wb_npc__T_8_data = 32'h0;
  assign queue_bits_wb_npc__T_8_addr = 6'h3;
  assign queue_bits_wb_npc__T_8_mask = 1'h0;
  assign queue_bits_wb_npc__T_8_en = 1'h0;
  assign queue_bits_wb_npc__T_9_data = 32'h0;
  assign queue_bits_wb_npc__T_9_addr = 6'h4;
  assign queue_bits_wb_npc__T_9_mask = 1'h0;
  assign queue_bits_wb_npc__T_9_en = 1'h0;
  assign queue_bits_wb_npc__T_10_data = 32'h0;
  assign queue_bits_wb_npc__T_10_addr = 6'h5;
  assign queue_bits_wb_npc__T_10_mask = 1'h0;
  assign queue_bits_wb_npc__T_10_en = 1'h0;
  assign queue_bits_wb_npc__T_11_data = 32'h0;
  assign queue_bits_wb_npc__T_11_addr = 6'h6;
  assign queue_bits_wb_npc__T_11_mask = 1'h0;
  assign queue_bits_wb_npc__T_11_en = 1'h0;
  assign queue_bits_wb_npc__T_12_data = 32'h0;
  assign queue_bits_wb_npc__T_12_addr = 6'h7;
  assign queue_bits_wb_npc__T_12_mask = 1'h0;
  assign queue_bits_wb_npc__T_12_en = 1'h0;
  assign queue_bits_wb_npc__T_13_data = 32'h0;
  assign queue_bits_wb_npc__T_13_addr = 6'h8;
  assign queue_bits_wb_npc__T_13_mask = 1'h0;
  assign queue_bits_wb_npc__T_13_en = 1'h0;
  assign queue_bits_wb_npc__T_14_data = 32'h0;
  assign queue_bits_wb_npc__T_14_addr = 6'h9;
  assign queue_bits_wb_npc__T_14_mask = 1'h0;
  assign queue_bits_wb_npc__T_14_en = 1'h0;
  assign queue_bits_wb_npc__T_15_data = 32'h0;
  assign queue_bits_wb_npc__T_15_addr = 6'ha;
  assign queue_bits_wb_npc__T_15_mask = 1'h0;
  assign queue_bits_wb_npc__T_15_en = 1'h0;
  assign queue_bits_wb_npc__T_16_data = 32'h0;
  assign queue_bits_wb_npc__T_16_addr = 6'hb;
  assign queue_bits_wb_npc__T_16_mask = 1'h0;
  assign queue_bits_wb_npc__T_16_en = 1'h0;
  assign queue_bits_wb_npc__T_17_data = 32'h0;
  assign queue_bits_wb_npc__T_17_addr = 6'hc;
  assign queue_bits_wb_npc__T_17_mask = 1'h0;
  assign queue_bits_wb_npc__T_17_en = 1'h0;
  assign queue_bits_wb_npc__T_18_data = 32'h0;
  assign queue_bits_wb_npc__T_18_addr = 6'hd;
  assign queue_bits_wb_npc__T_18_mask = 1'h0;
  assign queue_bits_wb_npc__T_18_en = 1'h0;
  assign queue_bits_wb_npc__T_19_data = 32'h0;
  assign queue_bits_wb_npc__T_19_addr = 6'he;
  assign queue_bits_wb_npc__T_19_mask = 1'h0;
  assign queue_bits_wb_npc__T_19_en = 1'h0;
  assign queue_bits_wb_npc__T_20_data = 32'h0;
  assign queue_bits_wb_npc__T_20_addr = 6'hf;
  assign queue_bits_wb_npc__T_20_mask = 1'h0;
  assign queue_bits_wb_npc__T_20_en = 1'h0;
  assign queue_bits_wb_npc__T_21_data = 32'h0;
  assign queue_bits_wb_npc__T_21_addr = 6'h10;
  assign queue_bits_wb_npc__T_21_mask = 1'h0;
  assign queue_bits_wb_npc__T_21_en = 1'h0;
  assign queue_bits_wb_npc__T_22_data = 32'h0;
  assign queue_bits_wb_npc__T_22_addr = 6'h11;
  assign queue_bits_wb_npc__T_22_mask = 1'h0;
  assign queue_bits_wb_npc__T_22_en = 1'h0;
  assign queue_bits_wb_npc__T_23_data = 32'h0;
  assign queue_bits_wb_npc__T_23_addr = 6'h12;
  assign queue_bits_wb_npc__T_23_mask = 1'h0;
  assign queue_bits_wb_npc__T_23_en = 1'h0;
  assign queue_bits_wb_npc__T_24_data = 32'h0;
  assign queue_bits_wb_npc__T_24_addr = 6'h13;
  assign queue_bits_wb_npc__T_24_mask = 1'h0;
  assign queue_bits_wb_npc__T_24_en = 1'h0;
  assign queue_bits_wb_npc__T_25_data = 32'h0;
  assign queue_bits_wb_npc__T_25_addr = 6'h14;
  assign queue_bits_wb_npc__T_25_mask = 1'h0;
  assign queue_bits_wb_npc__T_25_en = 1'h0;
  assign queue_bits_wb_npc__T_26_data = 32'h0;
  assign queue_bits_wb_npc__T_26_addr = 6'h15;
  assign queue_bits_wb_npc__T_26_mask = 1'h0;
  assign queue_bits_wb_npc__T_26_en = 1'h0;
  assign queue_bits_wb_npc__T_27_data = 32'h0;
  assign queue_bits_wb_npc__T_27_addr = 6'h16;
  assign queue_bits_wb_npc__T_27_mask = 1'h0;
  assign queue_bits_wb_npc__T_27_en = 1'h0;
  assign queue_bits_wb_npc__T_28_data = 32'h0;
  assign queue_bits_wb_npc__T_28_addr = 6'h17;
  assign queue_bits_wb_npc__T_28_mask = 1'h0;
  assign queue_bits_wb_npc__T_28_en = 1'h0;
  assign queue_bits_wb_npc__T_29_data = 32'h0;
  assign queue_bits_wb_npc__T_29_addr = 6'h18;
  assign queue_bits_wb_npc__T_29_mask = 1'h0;
  assign queue_bits_wb_npc__T_29_en = 1'h0;
  assign queue_bits_wb_npc__T_30_data = 32'h0;
  assign queue_bits_wb_npc__T_30_addr = 6'h19;
  assign queue_bits_wb_npc__T_30_mask = 1'h0;
  assign queue_bits_wb_npc__T_30_en = 1'h0;
  assign queue_bits_wb_npc__T_31_data = 32'h0;
  assign queue_bits_wb_npc__T_31_addr = 6'h1a;
  assign queue_bits_wb_npc__T_31_mask = 1'h0;
  assign queue_bits_wb_npc__T_31_en = 1'h0;
  assign queue_bits_wb_npc__T_32_data = 32'h0;
  assign queue_bits_wb_npc__T_32_addr = 6'h1b;
  assign queue_bits_wb_npc__T_32_mask = 1'h0;
  assign queue_bits_wb_npc__T_32_en = 1'h0;
  assign queue_bits_wb_npc__T_33_data = 32'h0;
  assign queue_bits_wb_npc__T_33_addr = 6'h1c;
  assign queue_bits_wb_npc__T_33_mask = 1'h0;
  assign queue_bits_wb_npc__T_33_en = 1'h0;
  assign queue_bits_wb_npc__T_34_data = 32'h0;
  assign queue_bits_wb_npc__T_34_addr = 6'h1d;
  assign queue_bits_wb_npc__T_34_mask = 1'h0;
  assign queue_bits_wb_npc__T_34_en = 1'h0;
  assign queue_bits_wb_npc__T_35_data = 32'h0;
  assign queue_bits_wb_npc__T_35_addr = 6'h1e;
  assign queue_bits_wb_npc__T_35_mask = 1'h0;
  assign queue_bits_wb_npc__T_35_en = 1'h0;
  assign queue_bits_wb_npc__T_36_data = 32'h0;
  assign queue_bits_wb_npc__T_36_addr = 6'h1f;
  assign queue_bits_wb_npc__T_36_mask = 1'h0;
  assign queue_bits_wb_npc__T_36_en = 1'h0;
  assign queue_bits_wb_npc__T_37_data = 32'h0;
  assign queue_bits_wb_npc__T_37_addr = 6'h20;
  assign queue_bits_wb_npc__T_37_mask = 1'h0;
  assign queue_bits_wb_npc__T_37_en = 1'h0;
  assign queue_bits_wb_npc__T_38_data = 32'h0;
  assign queue_bits_wb_npc__T_38_addr = 6'h21;
  assign queue_bits_wb_npc__T_38_mask = 1'h0;
  assign queue_bits_wb_npc__T_38_en = 1'h0;
  assign queue_bits_wb_npc__T_39_data = 32'h0;
  assign queue_bits_wb_npc__T_39_addr = 6'h22;
  assign queue_bits_wb_npc__T_39_mask = 1'h0;
  assign queue_bits_wb_npc__T_39_en = 1'h0;
  assign queue_bits_wb_npc__T_40_data = 32'h0;
  assign queue_bits_wb_npc__T_40_addr = 6'h23;
  assign queue_bits_wb_npc__T_40_mask = 1'h0;
  assign queue_bits_wb_npc__T_40_en = 1'h0;
  assign queue_bits_wb_npc__T_41_data = 32'h0;
  assign queue_bits_wb_npc__T_41_addr = 6'h24;
  assign queue_bits_wb_npc__T_41_mask = 1'h0;
  assign queue_bits_wb_npc__T_41_en = 1'h0;
  assign queue_bits_wb_npc__T_42_data = 32'h0;
  assign queue_bits_wb_npc__T_42_addr = 6'h25;
  assign queue_bits_wb_npc__T_42_mask = 1'h0;
  assign queue_bits_wb_npc__T_42_en = 1'h0;
  assign queue_bits_wb_npc__T_43_data = 32'h0;
  assign queue_bits_wb_npc__T_43_addr = 6'h26;
  assign queue_bits_wb_npc__T_43_mask = 1'h0;
  assign queue_bits_wb_npc__T_43_en = 1'h0;
  assign queue_bits_wb_npc__T_44_data = 32'h0;
  assign queue_bits_wb_npc__T_44_addr = 6'h27;
  assign queue_bits_wb_npc__T_44_mask = 1'h0;
  assign queue_bits_wb_npc__T_44_en = 1'h0;
  assign queue_bits_wb_npc__T_45_data = 32'h0;
  assign queue_bits_wb_npc__T_45_addr = 6'h28;
  assign queue_bits_wb_npc__T_45_mask = 1'h0;
  assign queue_bits_wb_npc__T_45_en = 1'h0;
  assign queue_bits_wb_npc__T_46_data = 32'h0;
  assign queue_bits_wb_npc__T_46_addr = 6'h29;
  assign queue_bits_wb_npc__T_46_mask = 1'h0;
  assign queue_bits_wb_npc__T_46_en = 1'h0;
  assign queue_bits_wb_npc__T_47_data = 32'h0;
  assign queue_bits_wb_npc__T_47_addr = 6'h2a;
  assign queue_bits_wb_npc__T_47_mask = 1'h0;
  assign queue_bits_wb_npc__T_47_en = 1'h0;
  assign queue_bits_wb_npc__T_48_data = 32'h0;
  assign queue_bits_wb_npc__T_48_addr = 6'h2b;
  assign queue_bits_wb_npc__T_48_mask = 1'h0;
  assign queue_bits_wb_npc__T_48_en = 1'h0;
  assign queue_bits_wb_npc__T_49_data = 32'h0;
  assign queue_bits_wb_npc__T_49_addr = 6'h2c;
  assign queue_bits_wb_npc__T_49_mask = 1'h0;
  assign queue_bits_wb_npc__T_49_en = 1'h0;
  assign queue_bits_wb_npc__T_50_data = 32'h0;
  assign queue_bits_wb_npc__T_50_addr = 6'h2d;
  assign queue_bits_wb_npc__T_50_mask = 1'h0;
  assign queue_bits_wb_npc__T_50_en = 1'h0;
  assign queue_bits_wb_npc__T_51_data = 32'h0;
  assign queue_bits_wb_npc__T_51_addr = 6'h2e;
  assign queue_bits_wb_npc__T_51_mask = 1'h0;
  assign queue_bits_wb_npc__T_51_en = 1'h0;
  assign queue_bits_wb_npc__T_52_data = 32'h0;
  assign queue_bits_wb_npc__T_52_addr = 6'h2f;
  assign queue_bits_wb_npc__T_52_mask = 1'h0;
  assign queue_bits_wb_npc__T_52_en = 1'h0;
  assign queue_bits_wb_npc__T_53_data = 32'h0;
  assign queue_bits_wb_npc__T_53_addr = 6'h30;
  assign queue_bits_wb_npc__T_53_mask = 1'h0;
  assign queue_bits_wb_npc__T_53_en = 1'h0;
  assign queue_bits_wb_npc__T_54_data = 32'h0;
  assign queue_bits_wb_npc__T_54_addr = 6'h31;
  assign queue_bits_wb_npc__T_54_mask = 1'h0;
  assign queue_bits_wb_npc__T_54_en = 1'h0;
  assign queue_bits_wb_npc__T_55_data = 32'h0;
  assign queue_bits_wb_npc__T_55_addr = 6'h32;
  assign queue_bits_wb_npc__T_55_mask = 1'h0;
  assign queue_bits_wb_npc__T_55_en = 1'h0;
  assign queue_bits_wb_npc__T_56_data = 32'h0;
  assign queue_bits_wb_npc__T_56_addr = 6'h33;
  assign queue_bits_wb_npc__T_56_mask = 1'h0;
  assign queue_bits_wb_npc__T_56_en = 1'h0;
  assign queue_bits_wb_npc__T_57_data = 32'h0;
  assign queue_bits_wb_npc__T_57_addr = 6'h34;
  assign queue_bits_wb_npc__T_57_mask = 1'h0;
  assign queue_bits_wb_npc__T_57_en = 1'h0;
  assign queue_bits_wb_npc__T_58_data = 32'h0;
  assign queue_bits_wb_npc__T_58_addr = 6'h35;
  assign queue_bits_wb_npc__T_58_mask = 1'h0;
  assign queue_bits_wb_npc__T_58_en = 1'h0;
  assign queue_bits_wb_npc__T_59_data = 32'h0;
  assign queue_bits_wb_npc__T_59_addr = 6'h36;
  assign queue_bits_wb_npc__T_59_mask = 1'h0;
  assign queue_bits_wb_npc__T_59_en = 1'h0;
  assign queue_bits_wb_npc__T_60_data = 32'h0;
  assign queue_bits_wb_npc__T_60_addr = 6'h37;
  assign queue_bits_wb_npc__T_60_mask = 1'h0;
  assign queue_bits_wb_npc__T_60_en = 1'h0;
  assign queue_bits_wb_npc__T_61_data = 32'h0;
  assign queue_bits_wb_npc__T_61_addr = 6'h38;
  assign queue_bits_wb_npc__T_61_mask = 1'h0;
  assign queue_bits_wb_npc__T_61_en = 1'h0;
  assign queue_bits_wb_npc__T_62_data = 32'h0;
  assign queue_bits_wb_npc__T_62_addr = 6'h39;
  assign queue_bits_wb_npc__T_62_mask = 1'h0;
  assign queue_bits_wb_npc__T_62_en = 1'h0;
  assign queue_bits_wb_npc__T_63_data = 32'h0;
  assign queue_bits_wb_npc__T_63_addr = 6'h3a;
  assign queue_bits_wb_npc__T_63_mask = 1'h0;
  assign queue_bits_wb_npc__T_63_en = 1'h0;
  assign queue_bits_wb_npc__T_64_data = 32'h0;
  assign queue_bits_wb_npc__T_64_addr = 6'h3b;
  assign queue_bits_wb_npc__T_64_mask = 1'h0;
  assign queue_bits_wb_npc__T_64_en = 1'h0;
  assign queue_bits_wb_npc__T_65_data = 32'h0;
  assign queue_bits_wb_npc__T_65_addr = 6'h3c;
  assign queue_bits_wb_npc__T_65_mask = 1'h0;
  assign queue_bits_wb_npc__T_65_en = 1'h0;
  assign queue_bits_wb_npc__T_66_data = 32'h0;
  assign queue_bits_wb_npc__T_66_addr = 6'h3d;
  assign queue_bits_wb_npc__T_66_mask = 1'h0;
  assign queue_bits_wb_npc__T_66_en = 1'h0;
  assign queue_bits_wb_npc__T_67_data = 32'h0;
  assign queue_bits_wb_npc__T_67_addr = 6'h3e;
  assign queue_bits_wb_npc__T_67_mask = 1'h0;
  assign queue_bits_wb_npc__T_67_en = 1'h0;
  assign queue_bits_wb_npc__T_68_data = 32'h0;
  assign queue_bits_wb_npc__T_68_addr = 6'h3f;
  assign queue_bits_wb_npc__T_68_mask = 1'h0;
  assign queue_bits_wb_npc__T_68_en = 1'h0;
  assign queue_bits_wb_npc__T_70_data = 32'h0;
  assign queue_bits_wb_npc__T_70_addr = 6'h0;
  assign queue_bits_wb_npc__T_70_mask = 1'h0;
  assign queue_bits_wb_npc__T_70_en = reset;
  assign queue_bits_wb_npc__T_71_data = 32'h0;
  assign queue_bits_wb_npc__T_71_addr = 6'h1;
  assign queue_bits_wb_npc__T_71_mask = 1'h0;
  assign queue_bits_wb_npc__T_71_en = reset;
  assign queue_bits_wb_npc__T_72_data = 32'h0;
  assign queue_bits_wb_npc__T_72_addr = 6'h2;
  assign queue_bits_wb_npc__T_72_mask = 1'h0;
  assign queue_bits_wb_npc__T_72_en = reset;
  assign queue_bits_wb_npc__T_73_data = 32'h0;
  assign queue_bits_wb_npc__T_73_addr = 6'h3;
  assign queue_bits_wb_npc__T_73_mask = 1'h0;
  assign queue_bits_wb_npc__T_73_en = reset;
  assign queue_bits_wb_npc__T_74_data = 32'h0;
  assign queue_bits_wb_npc__T_74_addr = 6'h4;
  assign queue_bits_wb_npc__T_74_mask = 1'h0;
  assign queue_bits_wb_npc__T_74_en = reset;
  assign queue_bits_wb_npc__T_75_data = 32'h0;
  assign queue_bits_wb_npc__T_75_addr = 6'h5;
  assign queue_bits_wb_npc__T_75_mask = 1'h0;
  assign queue_bits_wb_npc__T_75_en = reset;
  assign queue_bits_wb_npc__T_76_data = 32'h0;
  assign queue_bits_wb_npc__T_76_addr = 6'h6;
  assign queue_bits_wb_npc__T_76_mask = 1'h0;
  assign queue_bits_wb_npc__T_76_en = reset;
  assign queue_bits_wb_npc__T_77_data = 32'h0;
  assign queue_bits_wb_npc__T_77_addr = 6'h7;
  assign queue_bits_wb_npc__T_77_mask = 1'h0;
  assign queue_bits_wb_npc__T_77_en = reset;
  assign queue_bits_wb_npc__T_78_data = 32'h0;
  assign queue_bits_wb_npc__T_78_addr = 6'h8;
  assign queue_bits_wb_npc__T_78_mask = 1'h0;
  assign queue_bits_wb_npc__T_78_en = reset;
  assign queue_bits_wb_npc__T_79_data = 32'h0;
  assign queue_bits_wb_npc__T_79_addr = 6'h9;
  assign queue_bits_wb_npc__T_79_mask = 1'h0;
  assign queue_bits_wb_npc__T_79_en = reset;
  assign queue_bits_wb_npc__T_80_data = 32'h0;
  assign queue_bits_wb_npc__T_80_addr = 6'ha;
  assign queue_bits_wb_npc__T_80_mask = 1'h0;
  assign queue_bits_wb_npc__T_80_en = reset;
  assign queue_bits_wb_npc__T_81_data = 32'h0;
  assign queue_bits_wb_npc__T_81_addr = 6'hb;
  assign queue_bits_wb_npc__T_81_mask = 1'h0;
  assign queue_bits_wb_npc__T_81_en = reset;
  assign queue_bits_wb_npc__T_82_data = 32'h0;
  assign queue_bits_wb_npc__T_82_addr = 6'hc;
  assign queue_bits_wb_npc__T_82_mask = 1'h0;
  assign queue_bits_wb_npc__T_82_en = reset;
  assign queue_bits_wb_npc__T_83_data = 32'h0;
  assign queue_bits_wb_npc__T_83_addr = 6'hd;
  assign queue_bits_wb_npc__T_83_mask = 1'h0;
  assign queue_bits_wb_npc__T_83_en = reset;
  assign queue_bits_wb_npc__T_84_data = 32'h0;
  assign queue_bits_wb_npc__T_84_addr = 6'he;
  assign queue_bits_wb_npc__T_84_mask = 1'h0;
  assign queue_bits_wb_npc__T_84_en = reset;
  assign queue_bits_wb_npc__T_85_data = 32'h0;
  assign queue_bits_wb_npc__T_85_addr = 6'hf;
  assign queue_bits_wb_npc__T_85_mask = 1'h0;
  assign queue_bits_wb_npc__T_85_en = reset;
  assign queue_bits_wb_npc__T_86_data = 32'h0;
  assign queue_bits_wb_npc__T_86_addr = 6'h10;
  assign queue_bits_wb_npc__T_86_mask = 1'h0;
  assign queue_bits_wb_npc__T_86_en = reset;
  assign queue_bits_wb_npc__T_87_data = 32'h0;
  assign queue_bits_wb_npc__T_87_addr = 6'h11;
  assign queue_bits_wb_npc__T_87_mask = 1'h0;
  assign queue_bits_wb_npc__T_87_en = reset;
  assign queue_bits_wb_npc__T_88_data = 32'h0;
  assign queue_bits_wb_npc__T_88_addr = 6'h12;
  assign queue_bits_wb_npc__T_88_mask = 1'h0;
  assign queue_bits_wb_npc__T_88_en = reset;
  assign queue_bits_wb_npc__T_89_data = 32'h0;
  assign queue_bits_wb_npc__T_89_addr = 6'h13;
  assign queue_bits_wb_npc__T_89_mask = 1'h0;
  assign queue_bits_wb_npc__T_89_en = reset;
  assign queue_bits_wb_npc__T_90_data = 32'h0;
  assign queue_bits_wb_npc__T_90_addr = 6'h14;
  assign queue_bits_wb_npc__T_90_mask = 1'h0;
  assign queue_bits_wb_npc__T_90_en = reset;
  assign queue_bits_wb_npc__T_91_data = 32'h0;
  assign queue_bits_wb_npc__T_91_addr = 6'h15;
  assign queue_bits_wb_npc__T_91_mask = 1'h0;
  assign queue_bits_wb_npc__T_91_en = reset;
  assign queue_bits_wb_npc__T_92_data = 32'h0;
  assign queue_bits_wb_npc__T_92_addr = 6'h16;
  assign queue_bits_wb_npc__T_92_mask = 1'h0;
  assign queue_bits_wb_npc__T_92_en = reset;
  assign queue_bits_wb_npc__T_93_data = 32'h0;
  assign queue_bits_wb_npc__T_93_addr = 6'h17;
  assign queue_bits_wb_npc__T_93_mask = 1'h0;
  assign queue_bits_wb_npc__T_93_en = reset;
  assign queue_bits_wb_npc__T_94_data = 32'h0;
  assign queue_bits_wb_npc__T_94_addr = 6'h18;
  assign queue_bits_wb_npc__T_94_mask = 1'h0;
  assign queue_bits_wb_npc__T_94_en = reset;
  assign queue_bits_wb_npc__T_95_data = 32'h0;
  assign queue_bits_wb_npc__T_95_addr = 6'h19;
  assign queue_bits_wb_npc__T_95_mask = 1'h0;
  assign queue_bits_wb_npc__T_95_en = reset;
  assign queue_bits_wb_npc__T_96_data = 32'h0;
  assign queue_bits_wb_npc__T_96_addr = 6'h1a;
  assign queue_bits_wb_npc__T_96_mask = 1'h0;
  assign queue_bits_wb_npc__T_96_en = reset;
  assign queue_bits_wb_npc__T_97_data = 32'h0;
  assign queue_bits_wb_npc__T_97_addr = 6'h1b;
  assign queue_bits_wb_npc__T_97_mask = 1'h0;
  assign queue_bits_wb_npc__T_97_en = reset;
  assign queue_bits_wb_npc__T_98_data = 32'h0;
  assign queue_bits_wb_npc__T_98_addr = 6'h1c;
  assign queue_bits_wb_npc__T_98_mask = 1'h0;
  assign queue_bits_wb_npc__T_98_en = reset;
  assign queue_bits_wb_npc__T_99_data = 32'h0;
  assign queue_bits_wb_npc__T_99_addr = 6'h1d;
  assign queue_bits_wb_npc__T_99_mask = 1'h0;
  assign queue_bits_wb_npc__T_99_en = reset;
  assign queue_bits_wb_npc__T_100_data = 32'h0;
  assign queue_bits_wb_npc__T_100_addr = 6'h1e;
  assign queue_bits_wb_npc__T_100_mask = 1'h0;
  assign queue_bits_wb_npc__T_100_en = reset;
  assign queue_bits_wb_npc__T_101_data = 32'h0;
  assign queue_bits_wb_npc__T_101_addr = 6'h1f;
  assign queue_bits_wb_npc__T_101_mask = 1'h0;
  assign queue_bits_wb_npc__T_101_en = reset;
  assign queue_bits_wb_npc__T_102_data = 32'h0;
  assign queue_bits_wb_npc__T_102_addr = 6'h20;
  assign queue_bits_wb_npc__T_102_mask = 1'h0;
  assign queue_bits_wb_npc__T_102_en = reset;
  assign queue_bits_wb_npc__T_103_data = 32'h0;
  assign queue_bits_wb_npc__T_103_addr = 6'h21;
  assign queue_bits_wb_npc__T_103_mask = 1'h0;
  assign queue_bits_wb_npc__T_103_en = reset;
  assign queue_bits_wb_npc__T_104_data = 32'h0;
  assign queue_bits_wb_npc__T_104_addr = 6'h22;
  assign queue_bits_wb_npc__T_104_mask = 1'h0;
  assign queue_bits_wb_npc__T_104_en = reset;
  assign queue_bits_wb_npc__T_105_data = 32'h0;
  assign queue_bits_wb_npc__T_105_addr = 6'h23;
  assign queue_bits_wb_npc__T_105_mask = 1'h0;
  assign queue_bits_wb_npc__T_105_en = reset;
  assign queue_bits_wb_npc__T_106_data = 32'h0;
  assign queue_bits_wb_npc__T_106_addr = 6'h24;
  assign queue_bits_wb_npc__T_106_mask = 1'h0;
  assign queue_bits_wb_npc__T_106_en = reset;
  assign queue_bits_wb_npc__T_107_data = 32'h0;
  assign queue_bits_wb_npc__T_107_addr = 6'h25;
  assign queue_bits_wb_npc__T_107_mask = 1'h0;
  assign queue_bits_wb_npc__T_107_en = reset;
  assign queue_bits_wb_npc__T_108_data = 32'h0;
  assign queue_bits_wb_npc__T_108_addr = 6'h26;
  assign queue_bits_wb_npc__T_108_mask = 1'h0;
  assign queue_bits_wb_npc__T_108_en = reset;
  assign queue_bits_wb_npc__T_109_data = 32'h0;
  assign queue_bits_wb_npc__T_109_addr = 6'h27;
  assign queue_bits_wb_npc__T_109_mask = 1'h0;
  assign queue_bits_wb_npc__T_109_en = reset;
  assign queue_bits_wb_npc__T_110_data = 32'h0;
  assign queue_bits_wb_npc__T_110_addr = 6'h28;
  assign queue_bits_wb_npc__T_110_mask = 1'h0;
  assign queue_bits_wb_npc__T_110_en = reset;
  assign queue_bits_wb_npc__T_111_data = 32'h0;
  assign queue_bits_wb_npc__T_111_addr = 6'h29;
  assign queue_bits_wb_npc__T_111_mask = 1'h0;
  assign queue_bits_wb_npc__T_111_en = reset;
  assign queue_bits_wb_npc__T_112_data = 32'h0;
  assign queue_bits_wb_npc__T_112_addr = 6'h2a;
  assign queue_bits_wb_npc__T_112_mask = 1'h0;
  assign queue_bits_wb_npc__T_112_en = reset;
  assign queue_bits_wb_npc__T_113_data = 32'h0;
  assign queue_bits_wb_npc__T_113_addr = 6'h2b;
  assign queue_bits_wb_npc__T_113_mask = 1'h0;
  assign queue_bits_wb_npc__T_113_en = reset;
  assign queue_bits_wb_npc__T_114_data = 32'h0;
  assign queue_bits_wb_npc__T_114_addr = 6'h2c;
  assign queue_bits_wb_npc__T_114_mask = 1'h0;
  assign queue_bits_wb_npc__T_114_en = reset;
  assign queue_bits_wb_npc__T_115_data = 32'h0;
  assign queue_bits_wb_npc__T_115_addr = 6'h2d;
  assign queue_bits_wb_npc__T_115_mask = 1'h0;
  assign queue_bits_wb_npc__T_115_en = reset;
  assign queue_bits_wb_npc__T_116_data = 32'h0;
  assign queue_bits_wb_npc__T_116_addr = 6'h2e;
  assign queue_bits_wb_npc__T_116_mask = 1'h0;
  assign queue_bits_wb_npc__T_116_en = reset;
  assign queue_bits_wb_npc__T_117_data = 32'h0;
  assign queue_bits_wb_npc__T_117_addr = 6'h2f;
  assign queue_bits_wb_npc__T_117_mask = 1'h0;
  assign queue_bits_wb_npc__T_117_en = reset;
  assign queue_bits_wb_npc__T_118_data = 32'h0;
  assign queue_bits_wb_npc__T_118_addr = 6'h30;
  assign queue_bits_wb_npc__T_118_mask = 1'h0;
  assign queue_bits_wb_npc__T_118_en = reset;
  assign queue_bits_wb_npc__T_119_data = 32'h0;
  assign queue_bits_wb_npc__T_119_addr = 6'h31;
  assign queue_bits_wb_npc__T_119_mask = 1'h0;
  assign queue_bits_wb_npc__T_119_en = reset;
  assign queue_bits_wb_npc__T_120_data = 32'h0;
  assign queue_bits_wb_npc__T_120_addr = 6'h32;
  assign queue_bits_wb_npc__T_120_mask = 1'h0;
  assign queue_bits_wb_npc__T_120_en = reset;
  assign queue_bits_wb_npc__T_121_data = 32'h0;
  assign queue_bits_wb_npc__T_121_addr = 6'h33;
  assign queue_bits_wb_npc__T_121_mask = 1'h0;
  assign queue_bits_wb_npc__T_121_en = reset;
  assign queue_bits_wb_npc__T_122_data = 32'h0;
  assign queue_bits_wb_npc__T_122_addr = 6'h34;
  assign queue_bits_wb_npc__T_122_mask = 1'h0;
  assign queue_bits_wb_npc__T_122_en = reset;
  assign queue_bits_wb_npc__T_123_data = 32'h0;
  assign queue_bits_wb_npc__T_123_addr = 6'h35;
  assign queue_bits_wb_npc__T_123_mask = 1'h0;
  assign queue_bits_wb_npc__T_123_en = reset;
  assign queue_bits_wb_npc__T_124_data = 32'h0;
  assign queue_bits_wb_npc__T_124_addr = 6'h36;
  assign queue_bits_wb_npc__T_124_mask = 1'h0;
  assign queue_bits_wb_npc__T_124_en = reset;
  assign queue_bits_wb_npc__T_125_data = 32'h0;
  assign queue_bits_wb_npc__T_125_addr = 6'h37;
  assign queue_bits_wb_npc__T_125_mask = 1'h0;
  assign queue_bits_wb_npc__T_125_en = reset;
  assign queue_bits_wb_npc__T_126_data = 32'h0;
  assign queue_bits_wb_npc__T_126_addr = 6'h38;
  assign queue_bits_wb_npc__T_126_mask = 1'h0;
  assign queue_bits_wb_npc__T_126_en = reset;
  assign queue_bits_wb_npc__T_127_data = 32'h0;
  assign queue_bits_wb_npc__T_127_addr = 6'h39;
  assign queue_bits_wb_npc__T_127_mask = 1'h0;
  assign queue_bits_wb_npc__T_127_en = reset;
  assign queue_bits_wb_npc__T_128_data = 32'h0;
  assign queue_bits_wb_npc__T_128_addr = 6'h3a;
  assign queue_bits_wb_npc__T_128_mask = 1'h0;
  assign queue_bits_wb_npc__T_128_en = reset;
  assign queue_bits_wb_npc__T_129_data = 32'h0;
  assign queue_bits_wb_npc__T_129_addr = 6'h3b;
  assign queue_bits_wb_npc__T_129_mask = 1'h0;
  assign queue_bits_wb_npc__T_129_en = reset;
  assign queue_bits_wb_npc__T_130_data = 32'h0;
  assign queue_bits_wb_npc__T_130_addr = 6'h3c;
  assign queue_bits_wb_npc__T_130_mask = 1'h0;
  assign queue_bits_wb_npc__T_130_en = reset;
  assign queue_bits_wb_npc__T_131_data = 32'h0;
  assign queue_bits_wb_npc__T_131_addr = 6'h3d;
  assign queue_bits_wb_npc__T_131_mask = 1'h0;
  assign queue_bits_wb_npc__T_131_en = reset;
  assign queue_bits_wb_npc__T_132_data = 32'h0;
  assign queue_bits_wb_npc__T_132_addr = 6'h3e;
  assign queue_bits_wb_npc__T_132_mask = 1'h0;
  assign queue_bits_wb_npc__T_132_en = reset;
  assign queue_bits_wb_npc__T_133_data = 32'h0;
  assign queue_bits_wb_npc__T_133_addr = 6'h3f;
  assign queue_bits_wb_npc__T_133_mask = 1'h0;
  assign queue_bits_wb_npc__T_133_en = reset;
  assign queue_bits_wb_npc_q_head_w_data = 32'h0;
  assign queue_bits_wb_npc_q_head_w_addr = head;
  assign queue_bits_wb_npc_q_head_w_mask = 1'h0;
  assign queue_bits_wb_npc_q_head_w_en = io_deq_valid;
  assign io_deq_valid = queue_valid_q_head_r_data; // @[utils.scala 34:16]
  assign io_deq_bits_hi = queue_bits_hi_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_lo = queue_bits_lo_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_op1 = queue_bits_op1_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_fu_op = queue_bits_fu_op_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_id = queue_bits_wb_id_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_pc = queue_bits_wb_pc_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_instr_op = queue_bits_wb_instr_op_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_instr_rs_idx = queue_bits_wb_instr_rs_idx_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_instr_rt_idx = queue_bits_wb_instr_rt_idx_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_instr_rd_idx = queue_bits_wb_instr_rd_idx_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_instr_shamt = queue_bits_wb_instr_shamt_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_instr_func = queue_bits_wb_instr_func_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_rd_idx = queue_bits_wb_rd_idx_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_ip7 = queue_bits_wb_ip7_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_is_ds = queue_bits_wb_is_ds_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_is_br = queue_bits_wb_is_br_q_head_r_data; // @[utils.scala 35:15]
  assign io_deq_bits_wb_npc = queue_bits_wb_npc_q_head_r_data; // @[utils.scala 35:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_valid[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_hi[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_lo[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_op1[initvar] = _RAND_3[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_fu_op[initvar] = _RAND_4[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_id[initvar] = _RAND_5[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_pc[initvar] = _RAND_6[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_instr_op[initvar] = _RAND_7[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_instr_rs_idx[initvar] = _RAND_8[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_instr_rt_idx[initvar] = _RAND_9[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_10 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_instr_rd_idx[initvar] = _RAND_10[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_11 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_instr_shamt[initvar] = _RAND_11[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_instr_func[initvar] = _RAND_12[5:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_rd_idx[initvar] = _RAND_13[4:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_14 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_ip7[initvar] = _RAND_14[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_15 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_is_ds[initvar] = _RAND_15[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_is_br[initvar] = _RAND_16[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    queue_bits_wb_npc[initvar] = _RAND_17[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  head = _RAND_18[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(queue_valid__T_3_en & queue_valid__T_3_mask) begin
      queue_valid[queue_valid__T_3_addr] <= queue_valid__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_4_en & queue_valid__T_4_mask) begin
      queue_valid[queue_valid__T_4_addr] <= queue_valid__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_5_en & queue_valid__T_5_mask) begin
      queue_valid[queue_valid__T_5_addr] <= queue_valid__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_6_en & queue_valid__T_6_mask) begin
      queue_valid[queue_valid__T_6_addr] <= queue_valid__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_7_en & queue_valid__T_7_mask) begin
      queue_valid[queue_valid__T_7_addr] <= queue_valid__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_8_en & queue_valid__T_8_mask) begin
      queue_valid[queue_valid__T_8_addr] <= queue_valid__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_9_en & queue_valid__T_9_mask) begin
      queue_valid[queue_valid__T_9_addr] <= queue_valid__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_10_en & queue_valid__T_10_mask) begin
      queue_valid[queue_valid__T_10_addr] <= queue_valid__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_11_en & queue_valid__T_11_mask) begin
      queue_valid[queue_valid__T_11_addr] <= queue_valid__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_12_en & queue_valid__T_12_mask) begin
      queue_valid[queue_valid__T_12_addr] <= queue_valid__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_13_en & queue_valid__T_13_mask) begin
      queue_valid[queue_valid__T_13_addr] <= queue_valid__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_14_en & queue_valid__T_14_mask) begin
      queue_valid[queue_valid__T_14_addr] <= queue_valid__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_15_en & queue_valid__T_15_mask) begin
      queue_valid[queue_valid__T_15_addr] <= queue_valid__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_16_en & queue_valid__T_16_mask) begin
      queue_valid[queue_valid__T_16_addr] <= queue_valid__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_17_en & queue_valid__T_17_mask) begin
      queue_valid[queue_valid__T_17_addr] <= queue_valid__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_18_en & queue_valid__T_18_mask) begin
      queue_valid[queue_valid__T_18_addr] <= queue_valid__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_19_en & queue_valid__T_19_mask) begin
      queue_valid[queue_valid__T_19_addr] <= queue_valid__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_20_en & queue_valid__T_20_mask) begin
      queue_valid[queue_valid__T_20_addr] <= queue_valid__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_21_en & queue_valid__T_21_mask) begin
      queue_valid[queue_valid__T_21_addr] <= queue_valid__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_22_en & queue_valid__T_22_mask) begin
      queue_valid[queue_valid__T_22_addr] <= queue_valid__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_23_en & queue_valid__T_23_mask) begin
      queue_valid[queue_valid__T_23_addr] <= queue_valid__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_24_en & queue_valid__T_24_mask) begin
      queue_valid[queue_valid__T_24_addr] <= queue_valid__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_25_en & queue_valid__T_25_mask) begin
      queue_valid[queue_valid__T_25_addr] <= queue_valid__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_26_en & queue_valid__T_26_mask) begin
      queue_valid[queue_valid__T_26_addr] <= queue_valid__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_27_en & queue_valid__T_27_mask) begin
      queue_valid[queue_valid__T_27_addr] <= queue_valid__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_28_en & queue_valid__T_28_mask) begin
      queue_valid[queue_valid__T_28_addr] <= queue_valid__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_29_en & queue_valid__T_29_mask) begin
      queue_valid[queue_valid__T_29_addr] <= queue_valid__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_30_en & queue_valid__T_30_mask) begin
      queue_valid[queue_valid__T_30_addr] <= queue_valid__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_31_en & queue_valid__T_31_mask) begin
      queue_valid[queue_valid__T_31_addr] <= queue_valid__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_32_en & queue_valid__T_32_mask) begin
      queue_valid[queue_valid__T_32_addr] <= queue_valid__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_33_en & queue_valid__T_33_mask) begin
      queue_valid[queue_valid__T_33_addr] <= queue_valid__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_34_en & queue_valid__T_34_mask) begin
      queue_valid[queue_valid__T_34_addr] <= queue_valid__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_35_en & queue_valid__T_35_mask) begin
      queue_valid[queue_valid__T_35_addr] <= queue_valid__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_36_en & queue_valid__T_36_mask) begin
      queue_valid[queue_valid__T_36_addr] <= queue_valid__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_37_en & queue_valid__T_37_mask) begin
      queue_valid[queue_valid__T_37_addr] <= queue_valid__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_38_en & queue_valid__T_38_mask) begin
      queue_valid[queue_valid__T_38_addr] <= queue_valid__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_39_en & queue_valid__T_39_mask) begin
      queue_valid[queue_valid__T_39_addr] <= queue_valid__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_40_en & queue_valid__T_40_mask) begin
      queue_valid[queue_valid__T_40_addr] <= queue_valid__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_41_en & queue_valid__T_41_mask) begin
      queue_valid[queue_valid__T_41_addr] <= queue_valid__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_42_en & queue_valid__T_42_mask) begin
      queue_valid[queue_valid__T_42_addr] <= queue_valid__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_43_en & queue_valid__T_43_mask) begin
      queue_valid[queue_valid__T_43_addr] <= queue_valid__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_44_en & queue_valid__T_44_mask) begin
      queue_valid[queue_valid__T_44_addr] <= queue_valid__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_45_en & queue_valid__T_45_mask) begin
      queue_valid[queue_valid__T_45_addr] <= queue_valid__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_46_en & queue_valid__T_46_mask) begin
      queue_valid[queue_valid__T_46_addr] <= queue_valid__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_47_en & queue_valid__T_47_mask) begin
      queue_valid[queue_valid__T_47_addr] <= queue_valid__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_48_en & queue_valid__T_48_mask) begin
      queue_valid[queue_valid__T_48_addr] <= queue_valid__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_49_en & queue_valid__T_49_mask) begin
      queue_valid[queue_valid__T_49_addr] <= queue_valid__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_50_en & queue_valid__T_50_mask) begin
      queue_valid[queue_valid__T_50_addr] <= queue_valid__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_51_en & queue_valid__T_51_mask) begin
      queue_valid[queue_valid__T_51_addr] <= queue_valid__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_52_en & queue_valid__T_52_mask) begin
      queue_valid[queue_valid__T_52_addr] <= queue_valid__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_53_en & queue_valid__T_53_mask) begin
      queue_valid[queue_valid__T_53_addr] <= queue_valid__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_54_en & queue_valid__T_54_mask) begin
      queue_valid[queue_valid__T_54_addr] <= queue_valid__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_55_en & queue_valid__T_55_mask) begin
      queue_valid[queue_valid__T_55_addr] <= queue_valid__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_56_en & queue_valid__T_56_mask) begin
      queue_valid[queue_valid__T_56_addr] <= queue_valid__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_57_en & queue_valid__T_57_mask) begin
      queue_valid[queue_valid__T_57_addr] <= queue_valid__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_58_en & queue_valid__T_58_mask) begin
      queue_valid[queue_valid__T_58_addr] <= queue_valid__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_59_en & queue_valid__T_59_mask) begin
      queue_valid[queue_valid__T_59_addr] <= queue_valid__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_60_en & queue_valid__T_60_mask) begin
      queue_valid[queue_valid__T_60_addr] <= queue_valid__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_61_en & queue_valid__T_61_mask) begin
      queue_valid[queue_valid__T_61_addr] <= queue_valid__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_62_en & queue_valid__T_62_mask) begin
      queue_valid[queue_valid__T_62_addr] <= queue_valid__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_63_en & queue_valid__T_63_mask) begin
      queue_valid[queue_valid__T_63_addr] <= queue_valid__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_64_en & queue_valid__T_64_mask) begin
      queue_valid[queue_valid__T_64_addr] <= queue_valid__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_65_en & queue_valid__T_65_mask) begin
      queue_valid[queue_valid__T_65_addr] <= queue_valid__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_66_en & queue_valid__T_66_mask) begin
      queue_valid[queue_valid__T_66_addr] <= queue_valid__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_67_en & queue_valid__T_67_mask) begin
      queue_valid[queue_valid__T_67_addr] <= queue_valid__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_68_en & queue_valid__T_68_mask) begin
      queue_valid[queue_valid__T_68_addr] <= queue_valid__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_70_en & queue_valid__T_70_mask) begin
      queue_valid[queue_valid__T_70_addr] <= queue_valid__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_71_en & queue_valid__T_71_mask) begin
      queue_valid[queue_valid__T_71_addr] <= queue_valid__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_72_en & queue_valid__T_72_mask) begin
      queue_valid[queue_valid__T_72_addr] <= queue_valid__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_73_en & queue_valid__T_73_mask) begin
      queue_valid[queue_valid__T_73_addr] <= queue_valid__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_74_en & queue_valid__T_74_mask) begin
      queue_valid[queue_valid__T_74_addr] <= queue_valid__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_75_en & queue_valid__T_75_mask) begin
      queue_valid[queue_valid__T_75_addr] <= queue_valid__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_76_en & queue_valid__T_76_mask) begin
      queue_valid[queue_valid__T_76_addr] <= queue_valid__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_77_en & queue_valid__T_77_mask) begin
      queue_valid[queue_valid__T_77_addr] <= queue_valid__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_78_en & queue_valid__T_78_mask) begin
      queue_valid[queue_valid__T_78_addr] <= queue_valid__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_79_en & queue_valid__T_79_mask) begin
      queue_valid[queue_valid__T_79_addr] <= queue_valid__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_80_en & queue_valid__T_80_mask) begin
      queue_valid[queue_valid__T_80_addr] <= queue_valid__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_81_en & queue_valid__T_81_mask) begin
      queue_valid[queue_valid__T_81_addr] <= queue_valid__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_82_en & queue_valid__T_82_mask) begin
      queue_valid[queue_valid__T_82_addr] <= queue_valid__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_83_en & queue_valid__T_83_mask) begin
      queue_valid[queue_valid__T_83_addr] <= queue_valid__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_84_en & queue_valid__T_84_mask) begin
      queue_valid[queue_valid__T_84_addr] <= queue_valid__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_85_en & queue_valid__T_85_mask) begin
      queue_valid[queue_valid__T_85_addr] <= queue_valid__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_86_en & queue_valid__T_86_mask) begin
      queue_valid[queue_valid__T_86_addr] <= queue_valid__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_87_en & queue_valid__T_87_mask) begin
      queue_valid[queue_valid__T_87_addr] <= queue_valid__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_88_en & queue_valid__T_88_mask) begin
      queue_valid[queue_valid__T_88_addr] <= queue_valid__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_89_en & queue_valid__T_89_mask) begin
      queue_valid[queue_valid__T_89_addr] <= queue_valid__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_90_en & queue_valid__T_90_mask) begin
      queue_valid[queue_valid__T_90_addr] <= queue_valid__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_91_en & queue_valid__T_91_mask) begin
      queue_valid[queue_valid__T_91_addr] <= queue_valid__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_92_en & queue_valid__T_92_mask) begin
      queue_valid[queue_valid__T_92_addr] <= queue_valid__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_93_en & queue_valid__T_93_mask) begin
      queue_valid[queue_valid__T_93_addr] <= queue_valid__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_94_en & queue_valid__T_94_mask) begin
      queue_valid[queue_valid__T_94_addr] <= queue_valid__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_95_en & queue_valid__T_95_mask) begin
      queue_valid[queue_valid__T_95_addr] <= queue_valid__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_96_en & queue_valid__T_96_mask) begin
      queue_valid[queue_valid__T_96_addr] <= queue_valid__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_97_en & queue_valid__T_97_mask) begin
      queue_valid[queue_valid__T_97_addr] <= queue_valid__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_98_en & queue_valid__T_98_mask) begin
      queue_valid[queue_valid__T_98_addr] <= queue_valid__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_99_en & queue_valid__T_99_mask) begin
      queue_valid[queue_valid__T_99_addr] <= queue_valid__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_100_en & queue_valid__T_100_mask) begin
      queue_valid[queue_valid__T_100_addr] <= queue_valid__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_101_en & queue_valid__T_101_mask) begin
      queue_valid[queue_valid__T_101_addr] <= queue_valid__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_102_en & queue_valid__T_102_mask) begin
      queue_valid[queue_valid__T_102_addr] <= queue_valid__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_103_en & queue_valid__T_103_mask) begin
      queue_valid[queue_valid__T_103_addr] <= queue_valid__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_104_en & queue_valid__T_104_mask) begin
      queue_valid[queue_valid__T_104_addr] <= queue_valid__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_105_en & queue_valid__T_105_mask) begin
      queue_valid[queue_valid__T_105_addr] <= queue_valid__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_106_en & queue_valid__T_106_mask) begin
      queue_valid[queue_valid__T_106_addr] <= queue_valid__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_107_en & queue_valid__T_107_mask) begin
      queue_valid[queue_valid__T_107_addr] <= queue_valid__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_108_en & queue_valid__T_108_mask) begin
      queue_valid[queue_valid__T_108_addr] <= queue_valid__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_109_en & queue_valid__T_109_mask) begin
      queue_valid[queue_valid__T_109_addr] <= queue_valid__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_110_en & queue_valid__T_110_mask) begin
      queue_valid[queue_valid__T_110_addr] <= queue_valid__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_111_en & queue_valid__T_111_mask) begin
      queue_valid[queue_valid__T_111_addr] <= queue_valid__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_112_en & queue_valid__T_112_mask) begin
      queue_valid[queue_valid__T_112_addr] <= queue_valid__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_113_en & queue_valid__T_113_mask) begin
      queue_valid[queue_valid__T_113_addr] <= queue_valid__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_114_en & queue_valid__T_114_mask) begin
      queue_valid[queue_valid__T_114_addr] <= queue_valid__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_115_en & queue_valid__T_115_mask) begin
      queue_valid[queue_valid__T_115_addr] <= queue_valid__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_116_en & queue_valid__T_116_mask) begin
      queue_valid[queue_valid__T_116_addr] <= queue_valid__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_117_en & queue_valid__T_117_mask) begin
      queue_valid[queue_valid__T_117_addr] <= queue_valid__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_118_en & queue_valid__T_118_mask) begin
      queue_valid[queue_valid__T_118_addr] <= queue_valid__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_119_en & queue_valid__T_119_mask) begin
      queue_valid[queue_valid__T_119_addr] <= queue_valid__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_120_en & queue_valid__T_120_mask) begin
      queue_valid[queue_valid__T_120_addr] <= queue_valid__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_121_en & queue_valid__T_121_mask) begin
      queue_valid[queue_valid__T_121_addr] <= queue_valid__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_122_en & queue_valid__T_122_mask) begin
      queue_valid[queue_valid__T_122_addr] <= queue_valid__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_123_en & queue_valid__T_123_mask) begin
      queue_valid[queue_valid__T_123_addr] <= queue_valid__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_124_en & queue_valid__T_124_mask) begin
      queue_valid[queue_valid__T_124_addr] <= queue_valid__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_125_en & queue_valid__T_125_mask) begin
      queue_valid[queue_valid__T_125_addr] <= queue_valid__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_126_en & queue_valid__T_126_mask) begin
      queue_valid[queue_valid__T_126_addr] <= queue_valid__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_127_en & queue_valid__T_127_mask) begin
      queue_valid[queue_valid__T_127_addr] <= queue_valid__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_128_en & queue_valid__T_128_mask) begin
      queue_valid[queue_valid__T_128_addr] <= queue_valid__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_129_en & queue_valid__T_129_mask) begin
      queue_valid[queue_valid__T_129_addr] <= queue_valid__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_130_en & queue_valid__T_130_mask) begin
      queue_valid[queue_valid__T_130_addr] <= queue_valid__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_131_en & queue_valid__T_131_mask) begin
      queue_valid[queue_valid__T_131_addr] <= queue_valid__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_132_en & queue_valid__T_132_mask) begin
      queue_valid[queue_valid__T_132_addr] <= queue_valid__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_valid__T_133_en & queue_valid__T_133_mask) begin
      queue_valid[queue_valid__T_133_addr] <= queue_valid__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_valid_q_head_w_en & queue_valid_q_head_w_mask) begin
      queue_valid[queue_valid_q_head_w_addr] <= queue_valid_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_3_en & queue_bits_hi__T_3_mask) begin
      queue_bits_hi[queue_bits_hi__T_3_addr] <= queue_bits_hi__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_4_en & queue_bits_hi__T_4_mask) begin
      queue_bits_hi[queue_bits_hi__T_4_addr] <= queue_bits_hi__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_5_en & queue_bits_hi__T_5_mask) begin
      queue_bits_hi[queue_bits_hi__T_5_addr] <= queue_bits_hi__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_6_en & queue_bits_hi__T_6_mask) begin
      queue_bits_hi[queue_bits_hi__T_6_addr] <= queue_bits_hi__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_7_en & queue_bits_hi__T_7_mask) begin
      queue_bits_hi[queue_bits_hi__T_7_addr] <= queue_bits_hi__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_8_en & queue_bits_hi__T_8_mask) begin
      queue_bits_hi[queue_bits_hi__T_8_addr] <= queue_bits_hi__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_9_en & queue_bits_hi__T_9_mask) begin
      queue_bits_hi[queue_bits_hi__T_9_addr] <= queue_bits_hi__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_10_en & queue_bits_hi__T_10_mask) begin
      queue_bits_hi[queue_bits_hi__T_10_addr] <= queue_bits_hi__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_11_en & queue_bits_hi__T_11_mask) begin
      queue_bits_hi[queue_bits_hi__T_11_addr] <= queue_bits_hi__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_12_en & queue_bits_hi__T_12_mask) begin
      queue_bits_hi[queue_bits_hi__T_12_addr] <= queue_bits_hi__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_13_en & queue_bits_hi__T_13_mask) begin
      queue_bits_hi[queue_bits_hi__T_13_addr] <= queue_bits_hi__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_14_en & queue_bits_hi__T_14_mask) begin
      queue_bits_hi[queue_bits_hi__T_14_addr] <= queue_bits_hi__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_15_en & queue_bits_hi__T_15_mask) begin
      queue_bits_hi[queue_bits_hi__T_15_addr] <= queue_bits_hi__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_16_en & queue_bits_hi__T_16_mask) begin
      queue_bits_hi[queue_bits_hi__T_16_addr] <= queue_bits_hi__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_17_en & queue_bits_hi__T_17_mask) begin
      queue_bits_hi[queue_bits_hi__T_17_addr] <= queue_bits_hi__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_18_en & queue_bits_hi__T_18_mask) begin
      queue_bits_hi[queue_bits_hi__T_18_addr] <= queue_bits_hi__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_19_en & queue_bits_hi__T_19_mask) begin
      queue_bits_hi[queue_bits_hi__T_19_addr] <= queue_bits_hi__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_20_en & queue_bits_hi__T_20_mask) begin
      queue_bits_hi[queue_bits_hi__T_20_addr] <= queue_bits_hi__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_21_en & queue_bits_hi__T_21_mask) begin
      queue_bits_hi[queue_bits_hi__T_21_addr] <= queue_bits_hi__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_22_en & queue_bits_hi__T_22_mask) begin
      queue_bits_hi[queue_bits_hi__T_22_addr] <= queue_bits_hi__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_23_en & queue_bits_hi__T_23_mask) begin
      queue_bits_hi[queue_bits_hi__T_23_addr] <= queue_bits_hi__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_24_en & queue_bits_hi__T_24_mask) begin
      queue_bits_hi[queue_bits_hi__T_24_addr] <= queue_bits_hi__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_25_en & queue_bits_hi__T_25_mask) begin
      queue_bits_hi[queue_bits_hi__T_25_addr] <= queue_bits_hi__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_26_en & queue_bits_hi__T_26_mask) begin
      queue_bits_hi[queue_bits_hi__T_26_addr] <= queue_bits_hi__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_27_en & queue_bits_hi__T_27_mask) begin
      queue_bits_hi[queue_bits_hi__T_27_addr] <= queue_bits_hi__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_28_en & queue_bits_hi__T_28_mask) begin
      queue_bits_hi[queue_bits_hi__T_28_addr] <= queue_bits_hi__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_29_en & queue_bits_hi__T_29_mask) begin
      queue_bits_hi[queue_bits_hi__T_29_addr] <= queue_bits_hi__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_30_en & queue_bits_hi__T_30_mask) begin
      queue_bits_hi[queue_bits_hi__T_30_addr] <= queue_bits_hi__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_31_en & queue_bits_hi__T_31_mask) begin
      queue_bits_hi[queue_bits_hi__T_31_addr] <= queue_bits_hi__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_32_en & queue_bits_hi__T_32_mask) begin
      queue_bits_hi[queue_bits_hi__T_32_addr] <= queue_bits_hi__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_33_en & queue_bits_hi__T_33_mask) begin
      queue_bits_hi[queue_bits_hi__T_33_addr] <= queue_bits_hi__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_34_en & queue_bits_hi__T_34_mask) begin
      queue_bits_hi[queue_bits_hi__T_34_addr] <= queue_bits_hi__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_35_en & queue_bits_hi__T_35_mask) begin
      queue_bits_hi[queue_bits_hi__T_35_addr] <= queue_bits_hi__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_36_en & queue_bits_hi__T_36_mask) begin
      queue_bits_hi[queue_bits_hi__T_36_addr] <= queue_bits_hi__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_37_en & queue_bits_hi__T_37_mask) begin
      queue_bits_hi[queue_bits_hi__T_37_addr] <= queue_bits_hi__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_38_en & queue_bits_hi__T_38_mask) begin
      queue_bits_hi[queue_bits_hi__T_38_addr] <= queue_bits_hi__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_39_en & queue_bits_hi__T_39_mask) begin
      queue_bits_hi[queue_bits_hi__T_39_addr] <= queue_bits_hi__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_40_en & queue_bits_hi__T_40_mask) begin
      queue_bits_hi[queue_bits_hi__T_40_addr] <= queue_bits_hi__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_41_en & queue_bits_hi__T_41_mask) begin
      queue_bits_hi[queue_bits_hi__T_41_addr] <= queue_bits_hi__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_42_en & queue_bits_hi__T_42_mask) begin
      queue_bits_hi[queue_bits_hi__T_42_addr] <= queue_bits_hi__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_43_en & queue_bits_hi__T_43_mask) begin
      queue_bits_hi[queue_bits_hi__T_43_addr] <= queue_bits_hi__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_44_en & queue_bits_hi__T_44_mask) begin
      queue_bits_hi[queue_bits_hi__T_44_addr] <= queue_bits_hi__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_45_en & queue_bits_hi__T_45_mask) begin
      queue_bits_hi[queue_bits_hi__T_45_addr] <= queue_bits_hi__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_46_en & queue_bits_hi__T_46_mask) begin
      queue_bits_hi[queue_bits_hi__T_46_addr] <= queue_bits_hi__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_47_en & queue_bits_hi__T_47_mask) begin
      queue_bits_hi[queue_bits_hi__T_47_addr] <= queue_bits_hi__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_48_en & queue_bits_hi__T_48_mask) begin
      queue_bits_hi[queue_bits_hi__T_48_addr] <= queue_bits_hi__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_49_en & queue_bits_hi__T_49_mask) begin
      queue_bits_hi[queue_bits_hi__T_49_addr] <= queue_bits_hi__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_50_en & queue_bits_hi__T_50_mask) begin
      queue_bits_hi[queue_bits_hi__T_50_addr] <= queue_bits_hi__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_51_en & queue_bits_hi__T_51_mask) begin
      queue_bits_hi[queue_bits_hi__T_51_addr] <= queue_bits_hi__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_52_en & queue_bits_hi__T_52_mask) begin
      queue_bits_hi[queue_bits_hi__T_52_addr] <= queue_bits_hi__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_53_en & queue_bits_hi__T_53_mask) begin
      queue_bits_hi[queue_bits_hi__T_53_addr] <= queue_bits_hi__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_54_en & queue_bits_hi__T_54_mask) begin
      queue_bits_hi[queue_bits_hi__T_54_addr] <= queue_bits_hi__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_55_en & queue_bits_hi__T_55_mask) begin
      queue_bits_hi[queue_bits_hi__T_55_addr] <= queue_bits_hi__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_56_en & queue_bits_hi__T_56_mask) begin
      queue_bits_hi[queue_bits_hi__T_56_addr] <= queue_bits_hi__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_57_en & queue_bits_hi__T_57_mask) begin
      queue_bits_hi[queue_bits_hi__T_57_addr] <= queue_bits_hi__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_58_en & queue_bits_hi__T_58_mask) begin
      queue_bits_hi[queue_bits_hi__T_58_addr] <= queue_bits_hi__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_59_en & queue_bits_hi__T_59_mask) begin
      queue_bits_hi[queue_bits_hi__T_59_addr] <= queue_bits_hi__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_60_en & queue_bits_hi__T_60_mask) begin
      queue_bits_hi[queue_bits_hi__T_60_addr] <= queue_bits_hi__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_61_en & queue_bits_hi__T_61_mask) begin
      queue_bits_hi[queue_bits_hi__T_61_addr] <= queue_bits_hi__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_62_en & queue_bits_hi__T_62_mask) begin
      queue_bits_hi[queue_bits_hi__T_62_addr] <= queue_bits_hi__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_63_en & queue_bits_hi__T_63_mask) begin
      queue_bits_hi[queue_bits_hi__T_63_addr] <= queue_bits_hi__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_64_en & queue_bits_hi__T_64_mask) begin
      queue_bits_hi[queue_bits_hi__T_64_addr] <= queue_bits_hi__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_65_en & queue_bits_hi__T_65_mask) begin
      queue_bits_hi[queue_bits_hi__T_65_addr] <= queue_bits_hi__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_66_en & queue_bits_hi__T_66_mask) begin
      queue_bits_hi[queue_bits_hi__T_66_addr] <= queue_bits_hi__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_67_en & queue_bits_hi__T_67_mask) begin
      queue_bits_hi[queue_bits_hi__T_67_addr] <= queue_bits_hi__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_68_en & queue_bits_hi__T_68_mask) begin
      queue_bits_hi[queue_bits_hi__T_68_addr] <= queue_bits_hi__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_70_en & queue_bits_hi__T_70_mask) begin
      queue_bits_hi[queue_bits_hi__T_70_addr] <= queue_bits_hi__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_71_en & queue_bits_hi__T_71_mask) begin
      queue_bits_hi[queue_bits_hi__T_71_addr] <= queue_bits_hi__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_72_en & queue_bits_hi__T_72_mask) begin
      queue_bits_hi[queue_bits_hi__T_72_addr] <= queue_bits_hi__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_73_en & queue_bits_hi__T_73_mask) begin
      queue_bits_hi[queue_bits_hi__T_73_addr] <= queue_bits_hi__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_74_en & queue_bits_hi__T_74_mask) begin
      queue_bits_hi[queue_bits_hi__T_74_addr] <= queue_bits_hi__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_75_en & queue_bits_hi__T_75_mask) begin
      queue_bits_hi[queue_bits_hi__T_75_addr] <= queue_bits_hi__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_76_en & queue_bits_hi__T_76_mask) begin
      queue_bits_hi[queue_bits_hi__T_76_addr] <= queue_bits_hi__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_77_en & queue_bits_hi__T_77_mask) begin
      queue_bits_hi[queue_bits_hi__T_77_addr] <= queue_bits_hi__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_78_en & queue_bits_hi__T_78_mask) begin
      queue_bits_hi[queue_bits_hi__T_78_addr] <= queue_bits_hi__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_79_en & queue_bits_hi__T_79_mask) begin
      queue_bits_hi[queue_bits_hi__T_79_addr] <= queue_bits_hi__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_80_en & queue_bits_hi__T_80_mask) begin
      queue_bits_hi[queue_bits_hi__T_80_addr] <= queue_bits_hi__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_81_en & queue_bits_hi__T_81_mask) begin
      queue_bits_hi[queue_bits_hi__T_81_addr] <= queue_bits_hi__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_82_en & queue_bits_hi__T_82_mask) begin
      queue_bits_hi[queue_bits_hi__T_82_addr] <= queue_bits_hi__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_83_en & queue_bits_hi__T_83_mask) begin
      queue_bits_hi[queue_bits_hi__T_83_addr] <= queue_bits_hi__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_84_en & queue_bits_hi__T_84_mask) begin
      queue_bits_hi[queue_bits_hi__T_84_addr] <= queue_bits_hi__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_85_en & queue_bits_hi__T_85_mask) begin
      queue_bits_hi[queue_bits_hi__T_85_addr] <= queue_bits_hi__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_86_en & queue_bits_hi__T_86_mask) begin
      queue_bits_hi[queue_bits_hi__T_86_addr] <= queue_bits_hi__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_87_en & queue_bits_hi__T_87_mask) begin
      queue_bits_hi[queue_bits_hi__T_87_addr] <= queue_bits_hi__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_88_en & queue_bits_hi__T_88_mask) begin
      queue_bits_hi[queue_bits_hi__T_88_addr] <= queue_bits_hi__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_89_en & queue_bits_hi__T_89_mask) begin
      queue_bits_hi[queue_bits_hi__T_89_addr] <= queue_bits_hi__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_90_en & queue_bits_hi__T_90_mask) begin
      queue_bits_hi[queue_bits_hi__T_90_addr] <= queue_bits_hi__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_91_en & queue_bits_hi__T_91_mask) begin
      queue_bits_hi[queue_bits_hi__T_91_addr] <= queue_bits_hi__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_92_en & queue_bits_hi__T_92_mask) begin
      queue_bits_hi[queue_bits_hi__T_92_addr] <= queue_bits_hi__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_93_en & queue_bits_hi__T_93_mask) begin
      queue_bits_hi[queue_bits_hi__T_93_addr] <= queue_bits_hi__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_94_en & queue_bits_hi__T_94_mask) begin
      queue_bits_hi[queue_bits_hi__T_94_addr] <= queue_bits_hi__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_95_en & queue_bits_hi__T_95_mask) begin
      queue_bits_hi[queue_bits_hi__T_95_addr] <= queue_bits_hi__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_96_en & queue_bits_hi__T_96_mask) begin
      queue_bits_hi[queue_bits_hi__T_96_addr] <= queue_bits_hi__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_97_en & queue_bits_hi__T_97_mask) begin
      queue_bits_hi[queue_bits_hi__T_97_addr] <= queue_bits_hi__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_98_en & queue_bits_hi__T_98_mask) begin
      queue_bits_hi[queue_bits_hi__T_98_addr] <= queue_bits_hi__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_99_en & queue_bits_hi__T_99_mask) begin
      queue_bits_hi[queue_bits_hi__T_99_addr] <= queue_bits_hi__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_100_en & queue_bits_hi__T_100_mask) begin
      queue_bits_hi[queue_bits_hi__T_100_addr] <= queue_bits_hi__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_101_en & queue_bits_hi__T_101_mask) begin
      queue_bits_hi[queue_bits_hi__T_101_addr] <= queue_bits_hi__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_102_en & queue_bits_hi__T_102_mask) begin
      queue_bits_hi[queue_bits_hi__T_102_addr] <= queue_bits_hi__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_103_en & queue_bits_hi__T_103_mask) begin
      queue_bits_hi[queue_bits_hi__T_103_addr] <= queue_bits_hi__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_104_en & queue_bits_hi__T_104_mask) begin
      queue_bits_hi[queue_bits_hi__T_104_addr] <= queue_bits_hi__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_105_en & queue_bits_hi__T_105_mask) begin
      queue_bits_hi[queue_bits_hi__T_105_addr] <= queue_bits_hi__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_106_en & queue_bits_hi__T_106_mask) begin
      queue_bits_hi[queue_bits_hi__T_106_addr] <= queue_bits_hi__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_107_en & queue_bits_hi__T_107_mask) begin
      queue_bits_hi[queue_bits_hi__T_107_addr] <= queue_bits_hi__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_108_en & queue_bits_hi__T_108_mask) begin
      queue_bits_hi[queue_bits_hi__T_108_addr] <= queue_bits_hi__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_109_en & queue_bits_hi__T_109_mask) begin
      queue_bits_hi[queue_bits_hi__T_109_addr] <= queue_bits_hi__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_110_en & queue_bits_hi__T_110_mask) begin
      queue_bits_hi[queue_bits_hi__T_110_addr] <= queue_bits_hi__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_111_en & queue_bits_hi__T_111_mask) begin
      queue_bits_hi[queue_bits_hi__T_111_addr] <= queue_bits_hi__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_112_en & queue_bits_hi__T_112_mask) begin
      queue_bits_hi[queue_bits_hi__T_112_addr] <= queue_bits_hi__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_113_en & queue_bits_hi__T_113_mask) begin
      queue_bits_hi[queue_bits_hi__T_113_addr] <= queue_bits_hi__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_114_en & queue_bits_hi__T_114_mask) begin
      queue_bits_hi[queue_bits_hi__T_114_addr] <= queue_bits_hi__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_115_en & queue_bits_hi__T_115_mask) begin
      queue_bits_hi[queue_bits_hi__T_115_addr] <= queue_bits_hi__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_116_en & queue_bits_hi__T_116_mask) begin
      queue_bits_hi[queue_bits_hi__T_116_addr] <= queue_bits_hi__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_117_en & queue_bits_hi__T_117_mask) begin
      queue_bits_hi[queue_bits_hi__T_117_addr] <= queue_bits_hi__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_118_en & queue_bits_hi__T_118_mask) begin
      queue_bits_hi[queue_bits_hi__T_118_addr] <= queue_bits_hi__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_119_en & queue_bits_hi__T_119_mask) begin
      queue_bits_hi[queue_bits_hi__T_119_addr] <= queue_bits_hi__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_120_en & queue_bits_hi__T_120_mask) begin
      queue_bits_hi[queue_bits_hi__T_120_addr] <= queue_bits_hi__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_121_en & queue_bits_hi__T_121_mask) begin
      queue_bits_hi[queue_bits_hi__T_121_addr] <= queue_bits_hi__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_122_en & queue_bits_hi__T_122_mask) begin
      queue_bits_hi[queue_bits_hi__T_122_addr] <= queue_bits_hi__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_123_en & queue_bits_hi__T_123_mask) begin
      queue_bits_hi[queue_bits_hi__T_123_addr] <= queue_bits_hi__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_124_en & queue_bits_hi__T_124_mask) begin
      queue_bits_hi[queue_bits_hi__T_124_addr] <= queue_bits_hi__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_125_en & queue_bits_hi__T_125_mask) begin
      queue_bits_hi[queue_bits_hi__T_125_addr] <= queue_bits_hi__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_126_en & queue_bits_hi__T_126_mask) begin
      queue_bits_hi[queue_bits_hi__T_126_addr] <= queue_bits_hi__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_127_en & queue_bits_hi__T_127_mask) begin
      queue_bits_hi[queue_bits_hi__T_127_addr] <= queue_bits_hi__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_128_en & queue_bits_hi__T_128_mask) begin
      queue_bits_hi[queue_bits_hi__T_128_addr] <= queue_bits_hi__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_129_en & queue_bits_hi__T_129_mask) begin
      queue_bits_hi[queue_bits_hi__T_129_addr] <= queue_bits_hi__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_130_en & queue_bits_hi__T_130_mask) begin
      queue_bits_hi[queue_bits_hi__T_130_addr] <= queue_bits_hi__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_131_en & queue_bits_hi__T_131_mask) begin
      queue_bits_hi[queue_bits_hi__T_131_addr] <= queue_bits_hi__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_132_en & queue_bits_hi__T_132_mask) begin
      queue_bits_hi[queue_bits_hi__T_132_addr] <= queue_bits_hi__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi__T_133_en & queue_bits_hi__T_133_mask) begin
      queue_bits_hi[queue_bits_hi__T_133_addr] <= queue_bits_hi__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_hi_q_head_w_en & queue_bits_hi_q_head_w_mask) begin
      queue_bits_hi[queue_bits_hi_q_head_w_addr] <= queue_bits_hi_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_3_en & queue_bits_lo__T_3_mask) begin
      queue_bits_lo[queue_bits_lo__T_3_addr] <= queue_bits_lo__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_4_en & queue_bits_lo__T_4_mask) begin
      queue_bits_lo[queue_bits_lo__T_4_addr] <= queue_bits_lo__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_5_en & queue_bits_lo__T_5_mask) begin
      queue_bits_lo[queue_bits_lo__T_5_addr] <= queue_bits_lo__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_6_en & queue_bits_lo__T_6_mask) begin
      queue_bits_lo[queue_bits_lo__T_6_addr] <= queue_bits_lo__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_7_en & queue_bits_lo__T_7_mask) begin
      queue_bits_lo[queue_bits_lo__T_7_addr] <= queue_bits_lo__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_8_en & queue_bits_lo__T_8_mask) begin
      queue_bits_lo[queue_bits_lo__T_8_addr] <= queue_bits_lo__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_9_en & queue_bits_lo__T_9_mask) begin
      queue_bits_lo[queue_bits_lo__T_9_addr] <= queue_bits_lo__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_10_en & queue_bits_lo__T_10_mask) begin
      queue_bits_lo[queue_bits_lo__T_10_addr] <= queue_bits_lo__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_11_en & queue_bits_lo__T_11_mask) begin
      queue_bits_lo[queue_bits_lo__T_11_addr] <= queue_bits_lo__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_12_en & queue_bits_lo__T_12_mask) begin
      queue_bits_lo[queue_bits_lo__T_12_addr] <= queue_bits_lo__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_13_en & queue_bits_lo__T_13_mask) begin
      queue_bits_lo[queue_bits_lo__T_13_addr] <= queue_bits_lo__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_14_en & queue_bits_lo__T_14_mask) begin
      queue_bits_lo[queue_bits_lo__T_14_addr] <= queue_bits_lo__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_15_en & queue_bits_lo__T_15_mask) begin
      queue_bits_lo[queue_bits_lo__T_15_addr] <= queue_bits_lo__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_16_en & queue_bits_lo__T_16_mask) begin
      queue_bits_lo[queue_bits_lo__T_16_addr] <= queue_bits_lo__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_17_en & queue_bits_lo__T_17_mask) begin
      queue_bits_lo[queue_bits_lo__T_17_addr] <= queue_bits_lo__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_18_en & queue_bits_lo__T_18_mask) begin
      queue_bits_lo[queue_bits_lo__T_18_addr] <= queue_bits_lo__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_19_en & queue_bits_lo__T_19_mask) begin
      queue_bits_lo[queue_bits_lo__T_19_addr] <= queue_bits_lo__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_20_en & queue_bits_lo__T_20_mask) begin
      queue_bits_lo[queue_bits_lo__T_20_addr] <= queue_bits_lo__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_21_en & queue_bits_lo__T_21_mask) begin
      queue_bits_lo[queue_bits_lo__T_21_addr] <= queue_bits_lo__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_22_en & queue_bits_lo__T_22_mask) begin
      queue_bits_lo[queue_bits_lo__T_22_addr] <= queue_bits_lo__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_23_en & queue_bits_lo__T_23_mask) begin
      queue_bits_lo[queue_bits_lo__T_23_addr] <= queue_bits_lo__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_24_en & queue_bits_lo__T_24_mask) begin
      queue_bits_lo[queue_bits_lo__T_24_addr] <= queue_bits_lo__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_25_en & queue_bits_lo__T_25_mask) begin
      queue_bits_lo[queue_bits_lo__T_25_addr] <= queue_bits_lo__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_26_en & queue_bits_lo__T_26_mask) begin
      queue_bits_lo[queue_bits_lo__T_26_addr] <= queue_bits_lo__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_27_en & queue_bits_lo__T_27_mask) begin
      queue_bits_lo[queue_bits_lo__T_27_addr] <= queue_bits_lo__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_28_en & queue_bits_lo__T_28_mask) begin
      queue_bits_lo[queue_bits_lo__T_28_addr] <= queue_bits_lo__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_29_en & queue_bits_lo__T_29_mask) begin
      queue_bits_lo[queue_bits_lo__T_29_addr] <= queue_bits_lo__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_30_en & queue_bits_lo__T_30_mask) begin
      queue_bits_lo[queue_bits_lo__T_30_addr] <= queue_bits_lo__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_31_en & queue_bits_lo__T_31_mask) begin
      queue_bits_lo[queue_bits_lo__T_31_addr] <= queue_bits_lo__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_32_en & queue_bits_lo__T_32_mask) begin
      queue_bits_lo[queue_bits_lo__T_32_addr] <= queue_bits_lo__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_33_en & queue_bits_lo__T_33_mask) begin
      queue_bits_lo[queue_bits_lo__T_33_addr] <= queue_bits_lo__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_34_en & queue_bits_lo__T_34_mask) begin
      queue_bits_lo[queue_bits_lo__T_34_addr] <= queue_bits_lo__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_35_en & queue_bits_lo__T_35_mask) begin
      queue_bits_lo[queue_bits_lo__T_35_addr] <= queue_bits_lo__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_36_en & queue_bits_lo__T_36_mask) begin
      queue_bits_lo[queue_bits_lo__T_36_addr] <= queue_bits_lo__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_37_en & queue_bits_lo__T_37_mask) begin
      queue_bits_lo[queue_bits_lo__T_37_addr] <= queue_bits_lo__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_38_en & queue_bits_lo__T_38_mask) begin
      queue_bits_lo[queue_bits_lo__T_38_addr] <= queue_bits_lo__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_39_en & queue_bits_lo__T_39_mask) begin
      queue_bits_lo[queue_bits_lo__T_39_addr] <= queue_bits_lo__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_40_en & queue_bits_lo__T_40_mask) begin
      queue_bits_lo[queue_bits_lo__T_40_addr] <= queue_bits_lo__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_41_en & queue_bits_lo__T_41_mask) begin
      queue_bits_lo[queue_bits_lo__T_41_addr] <= queue_bits_lo__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_42_en & queue_bits_lo__T_42_mask) begin
      queue_bits_lo[queue_bits_lo__T_42_addr] <= queue_bits_lo__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_43_en & queue_bits_lo__T_43_mask) begin
      queue_bits_lo[queue_bits_lo__T_43_addr] <= queue_bits_lo__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_44_en & queue_bits_lo__T_44_mask) begin
      queue_bits_lo[queue_bits_lo__T_44_addr] <= queue_bits_lo__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_45_en & queue_bits_lo__T_45_mask) begin
      queue_bits_lo[queue_bits_lo__T_45_addr] <= queue_bits_lo__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_46_en & queue_bits_lo__T_46_mask) begin
      queue_bits_lo[queue_bits_lo__T_46_addr] <= queue_bits_lo__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_47_en & queue_bits_lo__T_47_mask) begin
      queue_bits_lo[queue_bits_lo__T_47_addr] <= queue_bits_lo__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_48_en & queue_bits_lo__T_48_mask) begin
      queue_bits_lo[queue_bits_lo__T_48_addr] <= queue_bits_lo__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_49_en & queue_bits_lo__T_49_mask) begin
      queue_bits_lo[queue_bits_lo__T_49_addr] <= queue_bits_lo__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_50_en & queue_bits_lo__T_50_mask) begin
      queue_bits_lo[queue_bits_lo__T_50_addr] <= queue_bits_lo__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_51_en & queue_bits_lo__T_51_mask) begin
      queue_bits_lo[queue_bits_lo__T_51_addr] <= queue_bits_lo__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_52_en & queue_bits_lo__T_52_mask) begin
      queue_bits_lo[queue_bits_lo__T_52_addr] <= queue_bits_lo__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_53_en & queue_bits_lo__T_53_mask) begin
      queue_bits_lo[queue_bits_lo__T_53_addr] <= queue_bits_lo__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_54_en & queue_bits_lo__T_54_mask) begin
      queue_bits_lo[queue_bits_lo__T_54_addr] <= queue_bits_lo__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_55_en & queue_bits_lo__T_55_mask) begin
      queue_bits_lo[queue_bits_lo__T_55_addr] <= queue_bits_lo__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_56_en & queue_bits_lo__T_56_mask) begin
      queue_bits_lo[queue_bits_lo__T_56_addr] <= queue_bits_lo__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_57_en & queue_bits_lo__T_57_mask) begin
      queue_bits_lo[queue_bits_lo__T_57_addr] <= queue_bits_lo__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_58_en & queue_bits_lo__T_58_mask) begin
      queue_bits_lo[queue_bits_lo__T_58_addr] <= queue_bits_lo__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_59_en & queue_bits_lo__T_59_mask) begin
      queue_bits_lo[queue_bits_lo__T_59_addr] <= queue_bits_lo__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_60_en & queue_bits_lo__T_60_mask) begin
      queue_bits_lo[queue_bits_lo__T_60_addr] <= queue_bits_lo__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_61_en & queue_bits_lo__T_61_mask) begin
      queue_bits_lo[queue_bits_lo__T_61_addr] <= queue_bits_lo__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_62_en & queue_bits_lo__T_62_mask) begin
      queue_bits_lo[queue_bits_lo__T_62_addr] <= queue_bits_lo__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_63_en & queue_bits_lo__T_63_mask) begin
      queue_bits_lo[queue_bits_lo__T_63_addr] <= queue_bits_lo__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_64_en & queue_bits_lo__T_64_mask) begin
      queue_bits_lo[queue_bits_lo__T_64_addr] <= queue_bits_lo__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_65_en & queue_bits_lo__T_65_mask) begin
      queue_bits_lo[queue_bits_lo__T_65_addr] <= queue_bits_lo__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_66_en & queue_bits_lo__T_66_mask) begin
      queue_bits_lo[queue_bits_lo__T_66_addr] <= queue_bits_lo__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_67_en & queue_bits_lo__T_67_mask) begin
      queue_bits_lo[queue_bits_lo__T_67_addr] <= queue_bits_lo__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_68_en & queue_bits_lo__T_68_mask) begin
      queue_bits_lo[queue_bits_lo__T_68_addr] <= queue_bits_lo__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_70_en & queue_bits_lo__T_70_mask) begin
      queue_bits_lo[queue_bits_lo__T_70_addr] <= queue_bits_lo__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_71_en & queue_bits_lo__T_71_mask) begin
      queue_bits_lo[queue_bits_lo__T_71_addr] <= queue_bits_lo__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_72_en & queue_bits_lo__T_72_mask) begin
      queue_bits_lo[queue_bits_lo__T_72_addr] <= queue_bits_lo__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_73_en & queue_bits_lo__T_73_mask) begin
      queue_bits_lo[queue_bits_lo__T_73_addr] <= queue_bits_lo__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_74_en & queue_bits_lo__T_74_mask) begin
      queue_bits_lo[queue_bits_lo__T_74_addr] <= queue_bits_lo__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_75_en & queue_bits_lo__T_75_mask) begin
      queue_bits_lo[queue_bits_lo__T_75_addr] <= queue_bits_lo__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_76_en & queue_bits_lo__T_76_mask) begin
      queue_bits_lo[queue_bits_lo__T_76_addr] <= queue_bits_lo__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_77_en & queue_bits_lo__T_77_mask) begin
      queue_bits_lo[queue_bits_lo__T_77_addr] <= queue_bits_lo__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_78_en & queue_bits_lo__T_78_mask) begin
      queue_bits_lo[queue_bits_lo__T_78_addr] <= queue_bits_lo__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_79_en & queue_bits_lo__T_79_mask) begin
      queue_bits_lo[queue_bits_lo__T_79_addr] <= queue_bits_lo__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_80_en & queue_bits_lo__T_80_mask) begin
      queue_bits_lo[queue_bits_lo__T_80_addr] <= queue_bits_lo__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_81_en & queue_bits_lo__T_81_mask) begin
      queue_bits_lo[queue_bits_lo__T_81_addr] <= queue_bits_lo__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_82_en & queue_bits_lo__T_82_mask) begin
      queue_bits_lo[queue_bits_lo__T_82_addr] <= queue_bits_lo__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_83_en & queue_bits_lo__T_83_mask) begin
      queue_bits_lo[queue_bits_lo__T_83_addr] <= queue_bits_lo__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_84_en & queue_bits_lo__T_84_mask) begin
      queue_bits_lo[queue_bits_lo__T_84_addr] <= queue_bits_lo__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_85_en & queue_bits_lo__T_85_mask) begin
      queue_bits_lo[queue_bits_lo__T_85_addr] <= queue_bits_lo__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_86_en & queue_bits_lo__T_86_mask) begin
      queue_bits_lo[queue_bits_lo__T_86_addr] <= queue_bits_lo__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_87_en & queue_bits_lo__T_87_mask) begin
      queue_bits_lo[queue_bits_lo__T_87_addr] <= queue_bits_lo__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_88_en & queue_bits_lo__T_88_mask) begin
      queue_bits_lo[queue_bits_lo__T_88_addr] <= queue_bits_lo__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_89_en & queue_bits_lo__T_89_mask) begin
      queue_bits_lo[queue_bits_lo__T_89_addr] <= queue_bits_lo__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_90_en & queue_bits_lo__T_90_mask) begin
      queue_bits_lo[queue_bits_lo__T_90_addr] <= queue_bits_lo__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_91_en & queue_bits_lo__T_91_mask) begin
      queue_bits_lo[queue_bits_lo__T_91_addr] <= queue_bits_lo__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_92_en & queue_bits_lo__T_92_mask) begin
      queue_bits_lo[queue_bits_lo__T_92_addr] <= queue_bits_lo__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_93_en & queue_bits_lo__T_93_mask) begin
      queue_bits_lo[queue_bits_lo__T_93_addr] <= queue_bits_lo__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_94_en & queue_bits_lo__T_94_mask) begin
      queue_bits_lo[queue_bits_lo__T_94_addr] <= queue_bits_lo__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_95_en & queue_bits_lo__T_95_mask) begin
      queue_bits_lo[queue_bits_lo__T_95_addr] <= queue_bits_lo__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_96_en & queue_bits_lo__T_96_mask) begin
      queue_bits_lo[queue_bits_lo__T_96_addr] <= queue_bits_lo__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_97_en & queue_bits_lo__T_97_mask) begin
      queue_bits_lo[queue_bits_lo__T_97_addr] <= queue_bits_lo__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_98_en & queue_bits_lo__T_98_mask) begin
      queue_bits_lo[queue_bits_lo__T_98_addr] <= queue_bits_lo__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_99_en & queue_bits_lo__T_99_mask) begin
      queue_bits_lo[queue_bits_lo__T_99_addr] <= queue_bits_lo__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_100_en & queue_bits_lo__T_100_mask) begin
      queue_bits_lo[queue_bits_lo__T_100_addr] <= queue_bits_lo__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_101_en & queue_bits_lo__T_101_mask) begin
      queue_bits_lo[queue_bits_lo__T_101_addr] <= queue_bits_lo__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_102_en & queue_bits_lo__T_102_mask) begin
      queue_bits_lo[queue_bits_lo__T_102_addr] <= queue_bits_lo__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_103_en & queue_bits_lo__T_103_mask) begin
      queue_bits_lo[queue_bits_lo__T_103_addr] <= queue_bits_lo__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_104_en & queue_bits_lo__T_104_mask) begin
      queue_bits_lo[queue_bits_lo__T_104_addr] <= queue_bits_lo__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_105_en & queue_bits_lo__T_105_mask) begin
      queue_bits_lo[queue_bits_lo__T_105_addr] <= queue_bits_lo__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_106_en & queue_bits_lo__T_106_mask) begin
      queue_bits_lo[queue_bits_lo__T_106_addr] <= queue_bits_lo__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_107_en & queue_bits_lo__T_107_mask) begin
      queue_bits_lo[queue_bits_lo__T_107_addr] <= queue_bits_lo__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_108_en & queue_bits_lo__T_108_mask) begin
      queue_bits_lo[queue_bits_lo__T_108_addr] <= queue_bits_lo__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_109_en & queue_bits_lo__T_109_mask) begin
      queue_bits_lo[queue_bits_lo__T_109_addr] <= queue_bits_lo__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_110_en & queue_bits_lo__T_110_mask) begin
      queue_bits_lo[queue_bits_lo__T_110_addr] <= queue_bits_lo__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_111_en & queue_bits_lo__T_111_mask) begin
      queue_bits_lo[queue_bits_lo__T_111_addr] <= queue_bits_lo__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_112_en & queue_bits_lo__T_112_mask) begin
      queue_bits_lo[queue_bits_lo__T_112_addr] <= queue_bits_lo__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_113_en & queue_bits_lo__T_113_mask) begin
      queue_bits_lo[queue_bits_lo__T_113_addr] <= queue_bits_lo__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_114_en & queue_bits_lo__T_114_mask) begin
      queue_bits_lo[queue_bits_lo__T_114_addr] <= queue_bits_lo__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_115_en & queue_bits_lo__T_115_mask) begin
      queue_bits_lo[queue_bits_lo__T_115_addr] <= queue_bits_lo__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_116_en & queue_bits_lo__T_116_mask) begin
      queue_bits_lo[queue_bits_lo__T_116_addr] <= queue_bits_lo__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_117_en & queue_bits_lo__T_117_mask) begin
      queue_bits_lo[queue_bits_lo__T_117_addr] <= queue_bits_lo__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_118_en & queue_bits_lo__T_118_mask) begin
      queue_bits_lo[queue_bits_lo__T_118_addr] <= queue_bits_lo__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_119_en & queue_bits_lo__T_119_mask) begin
      queue_bits_lo[queue_bits_lo__T_119_addr] <= queue_bits_lo__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_120_en & queue_bits_lo__T_120_mask) begin
      queue_bits_lo[queue_bits_lo__T_120_addr] <= queue_bits_lo__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_121_en & queue_bits_lo__T_121_mask) begin
      queue_bits_lo[queue_bits_lo__T_121_addr] <= queue_bits_lo__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_122_en & queue_bits_lo__T_122_mask) begin
      queue_bits_lo[queue_bits_lo__T_122_addr] <= queue_bits_lo__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_123_en & queue_bits_lo__T_123_mask) begin
      queue_bits_lo[queue_bits_lo__T_123_addr] <= queue_bits_lo__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_124_en & queue_bits_lo__T_124_mask) begin
      queue_bits_lo[queue_bits_lo__T_124_addr] <= queue_bits_lo__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_125_en & queue_bits_lo__T_125_mask) begin
      queue_bits_lo[queue_bits_lo__T_125_addr] <= queue_bits_lo__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_126_en & queue_bits_lo__T_126_mask) begin
      queue_bits_lo[queue_bits_lo__T_126_addr] <= queue_bits_lo__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_127_en & queue_bits_lo__T_127_mask) begin
      queue_bits_lo[queue_bits_lo__T_127_addr] <= queue_bits_lo__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_128_en & queue_bits_lo__T_128_mask) begin
      queue_bits_lo[queue_bits_lo__T_128_addr] <= queue_bits_lo__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_129_en & queue_bits_lo__T_129_mask) begin
      queue_bits_lo[queue_bits_lo__T_129_addr] <= queue_bits_lo__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_130_en & queue_bits_lo__T_130_mask) begin
      queue_bits_lo[queue_bits_lo__T_130_addr] <= queue_bits_lo__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_131_en & queue_bits_lo__T_131_mask) begin
      queue_bits_lo[queue_bits_lo__T_131_addr] <= queue_bits_lo__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_132_en & queue_bits_lo__T_132_mask) begin
      queue_bits_lo[queue_bits_lo__T_132_addr] <= queue_bits_lo__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo__T_133_en & queue_bits_lo__T_133_mask) begin
      queue_bits_lo[queue_bits_lo__T_133_addr] <= queue_bits_lo__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_lo_q_head_w_en & queue_bits_lo_q_head_w_mask) begin
      queue_bits_lo[queue_bits_lo_q_head_w_addr] <= queue_bits_lo_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_3_en & queue_bits_op1__T_3_mask) begin
      queue_bits_op1[queue_bits_op1__T_3_addr] <= queue_bits_op1__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_4_en & queue_bits_op1__T_4_mask) begin
      queue_bits_op1[queue_bits_op1__T_4_addr] <= queue_bits_op1__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_5_en & queue_bits_op1__T_5_mask) begin
      queue_bits_op1[queue_bits_op1__T_5_addr] <= queue_bits_op1__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_6_en & queue_bits_op1__T_6_mask) begin
      queue_bits_op1[queue_bits_op1__T_6_addr] <= queue_bits_op1__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_7_en & queue_bits_op1__T_7_mask) begin
      queue_bits_op1[queue_bits_op1__T_7_addr] <= queue_bits_op1__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_8_en & queue_bits_op1__T_8_mask) begin
      queue_bits_op1[queue_bits_op1__T_8_addr] <= queue_bits_op1__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_9_en & queue_bits_op1__T_9_mask) begin
      queue_bits_op1[queue_bits_op1__T_9_addr] <= queue_bits_op1__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_10_en & queue_bits_op1__T_10_mask) begin
      queue_bits_op1[queue_bits_op1__T_10_addr] <= queue_bits_op1__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_11_en & queue_bits_op1__T_11_mask) begin
      queue_bits_op1[queue_bits_op1__T_11_addr] <= queue_bits_op1__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_12_en & queue_bits_op1__T_12_mask) begin
      queue_bits_op1[queue_bits_op1__T_12_addr] <= queue_bits_op1__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_13_en & queue_bits_op1__T_13_mask) begin
      queue_bits_op1[queue_bits_op1__T_13_addr] <= queue_bits_op1__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_14_en & queue_bits_op1__T_14_mask) begin
      queue_bits_op1[queue_bits_op1__T_14_addr] <= queue_bits_op1__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_15_en & queue_bits_op1__T_15_mask) begin
      queue_bits_op1[queue_bits_op1__T_15_addr] <= queue_bits_op1__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_16_en & queue_bits_op1__T_16_mask) begin
      queue_bits_op1[queue_bits_op1__T_16_addr] <= queue_bits_op1__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_17_en & queue_bits_op1__T_17_mask) begin
      queue_bits_op1[queue_bits_op1__T_17_addr] <= queue_bits_op1__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_18_en & queue_bits_op1__T_18_mask) begin
      queue_bits_op1[queue_bits_op1__T_18_addr] <= queue_bits_op1__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_19_en & queue_bits_op1__T_19_mask) begin
      queue_bits_op1[queue_bits_op1__T_19_addr] <= queue_bits_op1__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_20_en & queue_bits_op1__T_20_mask) begin
      queue_bits_op1[queue_bits_op1__T_20_addr] <= queue_bits_op1__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_21_en & queue_bits_op1__T_21_mask) begin
      queue_bits_op1[queue_bits_op1__T_21_addr] <= queue_bits_op1__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_22_en & queue_bits_op1__T_22_mask) begin
      queue_bits_op1[queue_bits_op1__T_22_addr] <= queue_bits_op1__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_23_en & queue_bits_op1__T_23_mask) begin
      queue_bits_op1[queue_bits_op1__T_23_addr] <= queue_bits_op1__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_24_en & queue_bits_op1__T_24_mask) begin
      queue_bits_op1[queue_bits_op1__T_24_addr] <= queue_bits_op1__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_25_en & queue_bits_op1__T_25_mask) begin
      queue_bits_op1[queue_bits_op1__T_25_addr] <= queue_bits_op1__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_26_en & queue_bits_op1__T_26_mask) begin
      queue_bits_op1[queue_bits_op1__T_26_addr] <= queue_bits_op1__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_27_en & queue_bits_op1__T_27_mask) begin
      queue_bits_op1[queue_bits_op1__T_27_addr] <= queue_bits_op1__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_28_en & queue_bits_op1__T_28_mask) begin
      queue_bits_op1[queue_bits_op1__T_28_addr] <= queue_bits_op1__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_29_en & queue_bits_op1__T_29_mask) begin
      queue_bits_op1[queue_bits_op1__T_29_addr] <= queue_bits_op1__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_30_en & queue_bits_op1__T_30_mask) begin
      queue_bits_op1[queue_bits_op1__T_30_addr] <= queue_bits_op1__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_31_en & queue_bits_op1__T_31_mask) begin
      queue_bits_op1[queue_bits_op1__T_31_addr] <= queue_bits_op1__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_32_en & queue_bits_op1__T_32_mask) begin
      queue_bits_op1[queue_bits_op1__T_32_addr] <= queue_bits_op1__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_33_en & queue_bits_op1__T_33_mask) begin
      queue_bits_op1[queue_bits_op1__T_33_addr] <= queue_bits_op1__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_34_en & queue_bits_op1__T_34_mask) begin
      queue_bits_op1[queue_bits_op1__T_34_addr] <= queue_bits_op1__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_35_en & queue_bits_op1__T_35_mask) begin
      queue_bits_op1[queue_bits_op1__T_35_addr] <= queue_bits_op1__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_36_en & queue_bits_op1__T_36_mask) begin
      queue_bits_op1[queue_bits_op1__T_36_addr] <= queue_bits_op1__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_37_en & queue_bits_op1__T_37_mask) begin
      queue_bits_op1[queue_bits_op1__T_37_addr] <= queue_bits_op1__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_38_en & queue_bits_op1__T_38_mask) begin
      queue_bits_op1[queue_bits_op1__T_38_addr] <= queue_bits_op1__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_39_en & queue_bits_op1__T_39_mask) begin
      queue_bits_op1[queue_bits_op1__T_39_addr] <= queue_bits_op1__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_40_en & queue_bits_op1__T_40_mask) begin
      queue_bits_op1[queue_bits_op1__T_40_addr] <= queue_bits_op1__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_41_en & queue_bits_op1__T_41_mask) begin
      queue_bits_op1[queue_bits_op1__T_41_addr] <= queue_bits_op1__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_42_en & queue_bits_op1__T_42_mask) begin
      queue_bits_op1[queue_bits_op1__T_42_addr] <= queue_bits_op1__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_43_en & queue_bits_op1__T_43_mask) begin
      queue_bits_op1[queue_bits_op1__T_43_addr] <= queue_bits_op1__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_44_en & queue_bits_op1__T_44_mask) begin
      queue_bits_op1[queue_bits_op1__T_44_addr] <= queue_bits_op1__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_45_en & queue_bits_op1__T_45_mask) begin
      queue_bits_op1[queue_bits_op1__T_45_addr] <= queue_bits_op1__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_46_en & queue_bits_op1__T_46_mask) begin
      queue_bits_op1[queue_bits_op1__T_46_addr] <= queue_bits_op1__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_47_en & queue_bits_op1__T_47_mask) begin
      queue_bits_op1[queue_bits_op1__T_47_addr] <= queue_bits_op1__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_48_en & queue_bits_op1__T_48_mask) begin
      queue_bits_op1[queue_bits_op1__T_48_addr] <= queue_bits_op1__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_49_en & queue_bits_op1__T_49_mask) begin
      queue_bits_op1[queue_bits_op1__T_49_addr] <= queue_bits_op1__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_50_en & queue_bits_op1__T_50_mask) begin
      queue_bits_op1[queue_bits_op1__T_50_addr] <= queue_bits_op1__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_51_en & queue_bits_op1__T_51_mask) begin
      queue_bits_op1[queue_bits_op1__T_51_addr] <= queue_bits_op1__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_52_en & queue_bits_op1__T_52_mask) begin
      queue_bits_op1[queue_bits_op1__T_52_addr] <= queue_bits_op1__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_53_en & queue_bits_op1__T_53_mask) begin
      queue_bits_op1[queue_bits_op1__T_53_addr] <= queue_bits_op1__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_54_en & queue_bits_op1__T_54_mask) begin
      queue_bits_op1[queue_bits_op1__T_54_addr] <= queue_bits_op1__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_55_en & queue_bits_op1__T_55_mask) begin
      queue_bits_op1[queue_bits_op1__T_55_addr] <= queue_bits_op1__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_56_en & queue_bits_op1__T_56_mask) begin
      queue_bits_op1[queue_bits_op1__T_56_addr] <= queue_bits_op1__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_57_en & queue_bits_op1__T_57_mask) begin
      queue_bits_op1[queue_bits_op1__T_57_addr] <= queue_bits_op1__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_58_en & queue_bits_op1__T_58_mask) begin
      queue_bits_op1[queue_bits_op1__T_58_addr] <= queue_bits_op1__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_59_en & queue_bits_op1__T_59_mask) begin
      queue_bits_op1[queue_bits_op1__T_59_addr] <= queue_bits_op1__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_60_en & queue_bits_op1__T_60_mask) begin
      queue_bits_op1[queue_bits_op1__T_60_addr] <= queue_bits_op1__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_61_en & queue_bits_op1__T_61_mask) begin
      queue_bits_op1[queue_bits_op1__T_61_addr] <= queue_bits_op1__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_62_en & queue_bits_op1__T_62_mask) begin
      queue_bits_op1[queue_bits_op1__T_62_addr] <= queue_bits_op1__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_63_en & queue_bits_op1__T_63_mask) begin
      queue_bits_op1[queue_bits_op1__T_63_addr] <= queue_bits_op1__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_64_en & queue_bits_op1__T_64_mask) begin
      queue_bits_op1[queue_bits_op1__T_64_addr] <= queue_bits_op1__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_65_en & queue_bits_op1__T_65_mask) begin
      queue_bits_op1[queue_bits_op1__T_65_addr] <= queue_bits_op1__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_66_en & queue_bits_op1__T_66_mask) begin
      queue_bits_op1[queue_bits_op1__T_66_addr] <= queue_bits_op1__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_67_en & queue_bits_op1__T_67_mask) begin
      queue_bits_op1[queue_bits_op1__T_67_addr] <= queue_bits_op1__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_68_en & queue_bits_op1__T_68_mask) begin
      queue_bits_op1[queue_bits_op1__T_68_addr] <= queue_bits_op1__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_70_en & queue_bits_op1__T_70_mask) begin
      queue_bits_op1[queue_bits_op1__T_70_addr] <= queue_bits_op1__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_71_en & queue_bits_op1__T_71_mask) begin
      queue_bits_op1[queue_bits_op1__T_71_addr] <= queue_bits_op1__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_72_en & queue_bits_op1__T_72_mask) begin
      queue_bits_op1[queue_bits_op1__T_72_addr] <= queue_bits_op1__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_73_en & queue_bits_op1__T_73_mask) begin
      queue_bits_op1[queue_bits_op1__T_73_addr] <= queue_bits_op1__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_74_en & queue_bits_op1__T_74_mask) begin
      queue_bits_op1[queue_bits_op1__T_74_addr] <= queue_bits_op1__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_75_en & queue_bits_op1__T_75_mask) begin
      queue_bits_op1[queue_bits_op1__T_75_addr] <= queue_bits_op1__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_76_en & queue_bits_op1__T_76_mask) begin
      queue_bits_op1[queue_bits_op1__T_76_addr] <= queue_bits_op1__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_77_en & queue_bits_op1__T_77_mask) begin
      queue_bits_op1[queue_bits_op1__T_77_addr] <= queue_bits_op1__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_78_en & queue_bits_op1__T_78_mask) begin
      queue_bits_op1[queue_bits_op1__T_78_addr] <= queue_bits_op1__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_79_en & queue_bits_op1__T_79_mask) begin
      queue_bits_op1[queue_bits_op1__T_79_addr] <= queue_bits_op1__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_80_en & queue_bits_op1__T_80_mask) begin
      queue_bits_op1[queue_bits_op1__T_80_addr] <= queue_bits_op1__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_81_en & queue_bits_op1__T_81_mask) begin
      queue_bits_op1[queue_bits_op1__T_81_addr] <= queue_bits_op1__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_82_en & queue_bits_op1__T_82_mask) begin
      queue_bits_op1[queue_bits_op1__T_82_addr] <= queue_bits_op1__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_83_en & queue_bits_op1__T_83_mask) begin
      queue_bits_op1[queue_bits_op1__T_83_addr] <= queue_bits_op1__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_84_en & queue_bits_op1__T_84_mask) begin
      queue_bits_op1[queue_bits_op1__T_84_addr] <= queue_bits_op1__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_85_en & queue_bits_op1__T_85_mask) begin
      queue_bits_op1[queue_bits_op1__T_85_addr] <= queue_bits_op1__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_86_en & queue_bits_op1__T_86_mask) begin
      queue_bits_op1[queue_bits_op1__T_86_addr] <= queue_bits_op1__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_87_en & queue_bits_op1__T_87_mask) begin
      queue_bits_op1[queue_bits_op1__T_87_addr] <= queue_bits_op1__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_88_en & queue_bits_op1__T_88_mask) begin
      queue_bits_op1[queue_bits_op1__T_88_addr] <= queue_bits_op1__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_89_en & queue_bits_op1__T_89_mask) begin
      queue_bits_op1[queue_bits_op1__T_89_addr] <= queue_bits_op1__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_90_en & queue_bits_op1__T_90_mask) begin
      queue_bits_op1[queue_bits_op1__T_90_addr] <= queue_bits_op1__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_91_en & queue_bits_op1__T_91_mask) begin
      queue_bits_op1[queue_bits_op1__T_91_addr] <= queue_bits_op1__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_92_en & queue_bits_op1__T_92_mask) begin
      queue_bits_op1[queue_bits_op1__T_92_addr] <= queue_bits_op1__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_93_en & queue_bits_op1__T_93_mask) begin
      queue_bits_op1[queue_bits_op1__T_93_addr] <= queue_bits_op1__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_94_en & queue_bits_op1__T_94_mask) begin
      queue_bits_op1[queue_bits_op1__T_94_addr] <= queue_bits_op1__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_95_en & queue_bits_op1__T_95_mask) begin
      queue_bits_op1[queue_bits_op1__T_95_addr] <= queue_bits_op1__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_96_en & queue_bits_op1__T_96_mask) begin
      queue_bits_op1[queue_bits_op1__T_96_addr] <= queue_bits_op1__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_97_en & queue_bits_op1__T_97_mask) begin
      queue_bits_op1[queue_bits_op1__T_97_addr] <= queue_bits_op1__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_98_en & queue_bits_op1__T_98_mask) begin
      queue_bits_op1[queue_bits_op1__T_98_addr] <= queue_bits_op1__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_99_en & queue_bits_op1__T_99_mask) begin
      queue_bits_op1[queue_bits_op1__T_99_addr] <= queue_bits_op1__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_100_en & queue_bits_op1__T_100_mask) begin
      queue_bits_op1[queue_bits_op1__T_100_addr] <= queue_bits_op1__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_101_en & queue_bits_op1__T_101_mask) begin
      queue_bits_op1[queue_bits_op1__T_101_addr] <= queue_bits_op1__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_102_en & queue_bits_op1__T_102_mask) begin
      queue_bits_op1[queue_bits_op1__T_102_addr] <= queue_bits_op1__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_103_en & queue_bits_op1__T_103_mask) begin
      queue_bits_op1[queue_bits_op1__T_103_addr] <= queue_bits_op1__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_104_en & queue_bits_op1__T_104_mask) begin
      queue_bits_op1[queue_bits_op1__T_104_addr] <= queue_bits_op1__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_105_en & queue_bits_op1__T_105_mask) begin
      queue_bits_op1[queue_bits_op1__T_105_addr] <= queue_bits_op1__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_106_en & queue_bits_op1__T_106_mask) begin
      queue_bits_op1[queue_bits_op1__T_106_addr] <= queue_bits_op1__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_107_en & queue_bits_op1__T_107_mask) begin
      queue_bits_op1[queue_bits_op1__T_107_addr] <= queue_bits_op1__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_108_en & queue_bits_op1__T_108_mask) begin
      queue_bits_op1[queue_bits_op1__T_108_addr] <= queue_bits_op1__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_109_en & queue_bits_op1__T_109_mask) begin
      queue_bits_op1[queue_bits_op1__T_109_addr] <= queue_bits_op1__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_110_en & queue_bits_op1__T_110_mask) begin
      queue_bits_op1[queue_bits_op1__T_110_addr] <= queue_bits_op1__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_111_en & queue_bits_op1__T_111_mask) begin
      queue_bits_op1[queue_bits_op1__T_111_addr] <= queue_bits_op1__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_112_en & queue_bits_op1__T_112_mask) begin
      queue_bits_op1[queue_bits_op1__T_112_addr] <= queue_bits_op1__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_113_en & queue_bits_op1__T_113_mask) begin
      queue_bits_op1[queue_bits_op1__T_113_addr] <= queue_bits_op1__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_114_en & queue_bits_op1__T_114_mask) begin
      queue_bits_op1[queue_bits_op1__T_114_addr] <= queue_bits_op1__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_115_en & queue_bits_op1__T_115_mask) begin
      queue_bits_op1[queue_bits_op1__T_115_addr] <= queue_bits_op1__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_116_en & queue_bits_op1__T_116_mask) begin
      queue_bits_op1[queue_bits_op1__T_116_addr] <= queue_bits_op1__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_117_en & queue_bits_op1__T_117_mask) begin
      queue_bits_op1[queue_bits_op1__T_117_addr] <= queue_bits_op1__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_118_en & queue_bits_op1__T_118_mask) begin
      queue_bits_op1[queue_bits_op1__T_118_addr] <= queue_bits_op1__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_119_en & queue_bits_op1__T_119_mask) begin
      queue_bits_op1[queue_bits_op1__T_119_addr] <= queue_bits_op1__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_120_en & queue_bits_op1__T_120_mask) begin
      queue_bits_op1[queue_bits_op1__T_120_addr] <= queue_bits_op1__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_121_en & queue_bits_op1__T_121_mask) begin
      queue_bits_op1[queue_bits_op1__T_121_addr] <= queue_bits_op1__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_122_en & queue_bits_op1__T_122_mask) begin
      queue_bits_op1[queue_bits_op1__T_122_addr] <= queue_bits_op1__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_123_en & queue_bits_op1__T_123_mask) begin
      queue_bits_op1[queue_bits_op1__T_123_addr] <= queue_bits_op1__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_124_en & queue_bits_op1__T_124_mask) begin
      queue_bits_op1[queue_bits_op1__T_124_addr] <= queue_bits_op1__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_125_en & queue_bits_op1__T_125_mask) begin
      queue_bits_op1[queue_bits_op1__T_125_addr] <= queue_bits_op1__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_126_en & queue_bits_op1__T_126_mask) begin
      queue_bits_op1[queue_bits_op1__T_126_addr] <= queue_bits_op1__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_127_en & queue_bits_op1__T_127_mask) begin
      queue_bits_op1[queue_bits_op1__T_127_addr] <= queue_bits_op1__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_128_en & queue_bits_op1__T_128_mask) begin
      queue_bits_op1[queue_bits_op1__T_128_addr] <= queue_bits_op1__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_129_en & queue_bits_op1__T_129_mask) begin
      queue_bits_op1[queue_bits_op1__T_129_addr] <= queue_bits_op1__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_130_en & queue_bits_op1__T_130_mask) begin
      queue_bits_op1[queue_bits_op1__T_130_addr] <= queue_bits_op1__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_131_en & queue_bits_op1__T_131_mask) begin
      queue_bits_op1[queue_bits_op1__T_131_addr] <= queue_bits_op1__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_132_en & queue_bits_op1__T_132_mask) begin
      queue_bits_op1[queue_bits_op1__T_132_addr] <= queue_bits_op1__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1__T_133_en & queue_bits_op1__T_133_mask) begin
      queue_bits_op1[queue_bits_op1__T_133_addr] <= queue_bits_op1__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_op1_q_head_w_en & queue_bits_op1_q_head_w_mask) begin
      queue_bits_op1[queue_bits_op1_q_head_w_addr] <= queue_bits_op1_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_3_en & queue_bits_fu_op__T_3_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_3_addr] <= queue_bits_fu_op__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_4_en & queue_bits_fu_op__T_4_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_4_addr] <= queue_bits_fu_op__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_5_en & queue_bits_fu_op__T_5_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_5_addr] <= queue_bits_fu_op__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_6_en & queue_bits_fu_op__T_6_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_6_addr] <= queue_bits_fu_op__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_7_en & queue_bits_fu_op__T_7_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_7_addr] <= queue_bits_fu_op__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_8_en & queue_bits_fu_op__T_8_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_8_addr] <= queue_bits_fu_op__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_9_en & queue_bits_fu_op__T_9_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_9_addr] <= queue_bits_fu_op__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_10_en & queue_bits_fu_op__T_10_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_10_addr] <= queue_bits_fu_op__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_11_en & queue_bits_fu_op__T_11_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_11_addr] <= queue_bits_fu_op__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_12_en & queue_bits_fu_op__T_12_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_12_addr] <= queue_bits_fu_op__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_13_en & queue_bits_fu_op__T_13_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_13_addr] <= queue_bits_fu_op__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_14_en & queue_bits_fu_op__T_14_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_14_addr] <= queue_bits_fu_op__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_15_en & queue_bits_fu_op__T_15_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_15_addr] <= queue_bits_fu_op__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_16_en & queue_bits_fu_op__T_16_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_16_addr] <= queue_bits_fu_op__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_17_en & queue_bits_fu_op__T_17_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_17_addr] <= queue_bits_fu_op__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_18_en & queue_bits_fu_op__T_18_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_18_addr] <= queue_bits_fu_op__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_19_en & queue_bits_fu_op__T_19_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_19_addr] <= queue_bits_fu_op__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_20_en & queue_bits_fu_op__T_20_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_20_addr] <= queue_bits_fu_op__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_21_en & queue_bits_fu_op__T_21_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_21_addr] <= queue_bits_fu_op__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_22_en & queue_bits_fu_op__T_22_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_22_addr] <= queue_bits_fu_op__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_23_en & queue_bits_fu_op__T_23_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_23_addr] <= queue_bits_fu_op__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_24_en & queue_bits_fu_op__T_24_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_24_addr] <= queue_bits_fu_op__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_25_en & queue_bits_fu_op__T_25_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_25_addr] <= queue_bits_fu_op__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_26_en & queue_bits_fu_op__T_26_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_26_addr] <= queue_bits_fu_op__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_27_en & queue_bits_fu_op__T_27_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_27_addr] <= queue_bits_fu_op__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_28_en & queue_bits_fu_op__T_28_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_28_addr] <= queue_bits_fu_op__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_29_en & queue_bits_fu_op__T_29_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_29_addr] <= queue_bits_fu_op__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_30_en & queue_bits_fu_op__T_30_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_30_addr] <= queue_bits_fu_op__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_31_en & queue_bits_fu_op__T_31_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_31_addr] <= queue_bits_fu_op__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_32_en & queue_bits_fu_op__T_32_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_32_addr] <= queue_bits_fu_op__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_33_en & queue_bits_fu_op__T_33_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_33_addr] <= queue_bits_fu_op__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_34_en & queue_bits_fu_op__T_34_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_34_addr] <= queue_bits_fu_op__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_35_en & queue_bits_fu_op__T_35_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_35_addr] <= queue_bits_fu_op__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_36_en & queue_bits_fu_op__T_36_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_36_addr] <= queue_bits_fu_op__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_37_en & queue_bits_fu_op__T_37_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_37_addr] <= queue_bits_fu_op__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_38_en & queue_bits_fu_op__T_38_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_38_addr] <= queue_bits_fu_op__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_39_en & queue_bits_fu_op__T_39_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_39_addr] <= queue_bits_fu_op__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_40_en & queue_bits_fu_op__T_40_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_40_addr] <= queue_bits_fu_op__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_41_en & queue_bits_fu_op__T_41_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_41_addr] <= queue_bits_fu_op__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_42_en & queue_bits_fu_op__T_42_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_42_addr] <= queue_bits_fu_op__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_43_en & queue_bits_fu_op__T_43_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_43_addr] <= queue_bits_fu_op__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_44_en & queue_bits_fu_op__T_44_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_44_addr] <= queue_bits_fu_op__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_45_en & queue_bits_fu_op__T_45_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_45_addr] <= queue_bits_fu_op__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_46_en & queue_bits_fu_op__T_46_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_46_addr] <= queue_bits_fu_op__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_47_en & queue_bits_fu_op__T_47_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_47_addr] <= queue_bits_fu_op__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_48_en & queue_bits_fu_op__T_48_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_48_addr] <= queue_bits_fu_op__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_49_en & queue_bits_fu_op__T_49_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_49_addr] <= queue_bits_fu_op__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_50_en & queue_bits_fu_op__T_50_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_50_addr] <= queue_bits_fu_op__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_51_en & queue_bits_fu_op__T_51_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_51_addr] <= queue_bits_fu_op__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_52_en & queue_bits_fu_op__T_52_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_52_addr] <= queue_bits_fu_op__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_53_en & queue_bits_fu_op__T_53_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_53_addr] <= queue_bits_fu_op__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_54_en & queue_bits_fu_op__T_54_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_54_addr] <= queue_bits_fu_op__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_55_en & queue_bits_fu_op__T_55_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_55_addr] <= queue_bits_fu_op__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_56_en & queue_bits_fu_op__T_56_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_56_addr] <= queue_bits_fu_op__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_57_en & queue_bits_fu_op__T_57_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_57_addr] <= queue_bits_fu_op__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_58_en & queue_bits_fu_op__T_58_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_58_addr] <= queue_bits_fu_op__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_59_en & queue_bits_fu_op__T_59_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_59_addr] <= queue_bits_fu_op__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_60_en & queue_bits_fu_op__T_60_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_60_addr] <= queue_bits_fu_op__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_61_en & queue_bits_fu_op__T_61_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_61_addr] <= queue_bits_fu_op__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_62_en & queue_bits_fu_op__T_62_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_62_addr] <= queue_bits_fu_op__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_63_en & queue_bits_fu_op__T_63_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_63_addr] <= queue_bits_fu_op__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_64_en & queue_bits_fu_op__T_64_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_64_addr] <= queue_bits_fu_op__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_65_en & queue_bits_fu_op__T_65_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_65_addr] <= queue_bits_fu_op__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_66_en & queue_bits_fu_op__T_66_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_66_addr] <= queue_bits_fu_op__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_67_en & queue_bits_fu_op__T_67_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_67_addr] <= queue_bits_fu_op__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_68_en & queue_bits_fu_op__T_68_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_68_addr] <= queue_bits_fu_op__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_70_en & queue_bits_fu_op__T_70_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_70_addr] <= queue_bits_fu_op__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_71_en & queue_bits_fu_op__T_71_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_71_addr] <= queue_bits_fu_op__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_72_en & queue_bits_fu_op__T_72_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_72_addr] <= queue_bits_fu_op__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_73_en & queue_bits_fu_op__T_73_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_73_addr] <= queue_bits_fu_op__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_74_en & queue_bits_fu_op__T_74_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_74_addr] <= queue_bits_fu_op__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_75_en & queue_bits_fu_op__T_75_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_75_addr] <= queue_bits_fu_op__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_76_en & queue_bits_fu_op__T_76_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_76_addr] <= queue_bits_fu_op__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_77_en & queue_bits_fu_op__T_77_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_77_addr] <= queue_bits_fu_op__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_78_en & queue_bits_fu_op__T_78_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_78_addr] <= queue_bits_fu_op__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_79_en & queue_bits_fu_op__T_79_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_79_addr] <= queue_bits_fu_op__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_80_en & queue_bits_fu_op__T_80_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_80_addr] <= queue_bits_fu_op__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_81_en & queue_bits_fu_op__T_81_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_81_addr] <= queue_bits_fu_op__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_82_en & queue_bits_fu_op__T_82_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_82_addr] <= queue_bits_fu_op__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_83_en & queue_bits_fu_op__T_83_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_83_addr] <= queue_bits_fu_op__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_84_en & queue_bits_fu_op__T_84_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_84_addr] <= queue_bits_fu_op__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_85_en & queue_bits_fu_op__T_85_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_85_addr] <= queue_bits_fu_op__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_86_en & queue_bits_fu_op__T_86_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_86_addr] <= queue_bits_fu_op__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_87_en & queue_bits_fu_op__T_87_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_87_addr] <= queue_bits_fu_op__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_88_en & queue_bits_fu_op__T_88_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_88_addr] <= queue_bits_fu_op__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_89_en & queue_bits_fu_op__T_89_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_89_addr] <= queue_bits_fu_op__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_90_en & queue_bits_fu_op__T_90_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_90_addr] <= queue_bits_fu_op__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_91_en & queue_bits_fu_op__T_91_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_91_addr] <= queue_bits_fu_op__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_92_en & queue_bits_fu_op__T_92_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_92_addr] <= queue_bits_fu_op__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_93_en & queue_bits_fu_op__T_93_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_93_addr] <= queue_bits_fu_op__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_94_en & queue_bits_fu_op__T_94_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_94_addr] <= queue_bits_fu_op__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_95_en & queue_bits_fu_op__T_95_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_95_addr] <= queue_bits_fu_op__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_96_en & queue_bits_fu_op__T_96_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_96_addr] <= queue_bits_fu_op__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_97_en & queue_bits_fu_op__T_97_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_97_addr] <= queue_bits_fu_op__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_98_en & queue_bits_fu_op__T_98_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_98_addr] <= queue_bits_fu_op__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_99_en & queue_bits_fu_op__T_99_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_99_addr] <= queue_bits_fu_op__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_100_en & queue_bits_fu_op__T_100_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_100_addr] <= queue_bits_fu_op__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_101_en & queue_bits_fu_op__T_101_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_101_addr] <= queue_bits_fu_op__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_102_en & queue_bits_fu_op__T_102_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_102_addr] <= queue_bits_fu_op__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_103_en & queue_bits_fu_op__T_103_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_103_addr] <= queue_bits_fu_op__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_104_en & queue_bits_fu_op__T_104_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_104_addr] <= queue_bits_fu_op__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_105_en & queue_bits_fu_op__T_105_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_105_addr] <= queue_bits_fu_op__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_106_en & queue_bits_fu_op__T_106_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_106_addr] <= queue_bits_fu_op__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_107_en & queue_bits_fu_op__T_107_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_107_addr] <= queue_bits_fu_op__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_108_en & queue_bits_fu_op__T_108_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_108_addr] <= queue_bits_fu_op__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_109_en & queue_bits_fu_op__T_109_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_109_addr] <= queue_bits_fu_op__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_110_en & queue_bits_fu_op__T_110_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_110_addr] <= queue_bits_fu_op__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_111_en & queue_bits_fu_op__T_111_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_111_addr] <= queue_bits_fu_op__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_112_en & queue_bits_fu_op__T_112_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_112_addr] <= queue_bits_fu_op__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_113_en & queue_bits_fu_op__T_113_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_113_addr] <= queue_bits_fu_op__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_114_en & queue_bits_fu_op__T_114_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_114_addr] <= queue_bits_fu_op__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_115_en & queue_bits_fu_op__T_115_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_115_addr] <= queue_bits_fu_op__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_116_en & queue_bits_fu_op__T_116_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_116_addr] <= queue_bits_fu_op__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_117_en & queue_bits_fu_op__T_117_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_117_addr] <= queue_bits_fu_op__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_118_en & queue_bits_fu_op__T_118_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_118_addr] <= queue_bits_fu_op__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_119_en & queue_bits_fu_op__T_119_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_119_addr] <= queue_bits_fu_op__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_120_en & queue_bits_fu_op__T_120_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_120_addr] <= queue_bits_fu_op__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_121_en & queue_bits_fu_op__T_121_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_121_addr] <= queue_bits_fu_op__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_122_en & queue_bits_fu_op__T_122_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_122_addr] <= queue_bits_fu_op__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_123_en & queue_bits_fu_op__T_123_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_123_addr] <= queue_bits_fu_op__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_124_en & queue_bits_fu_op__T_124_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_124_addr] <= queue_bits_fu_op__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_125_en & queue_bits_fu_op__T_125_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_125_addr] <= queue_bits_fu_op__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_126_en & queue_bits_fu_op__T_126_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_126_addr] <= queue_bits_fu_op__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_127_en & queue_bits_fu_op__T_127_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_127_addr] <= queue_bits_fu_op__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_128_en & queue_bits_fu_op__T_128_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_128_addr] <= queue_bits_fu_op__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_129_en & queue_bits_fu_op__T_129_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_129_addr] <= queue_bits_fu_op__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_130_en & queue_bits_fu_op__T_130_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_130_addr] <= queue_bits_fu_op__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_131_en & queue_bits_fu_op__T_131_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_131_addr] <= queue_bits_fu_op__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_132_en & queue_bits_fu_op__T_132_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_132_addr] <= queue_bits_fu_op__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op__T_133_en & queue_bits_fu_op__T_133_mask) begin
      queue_bits_fu_op[queue_bits_fu_op__T_133_addr] <= queue_bits_fu_op__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_fu_op_q_head_w_en & queue_bits_fu_op_q_head_w_mask) begin
      queue_bits_fu_op[queue_bits_fu_op_q_head_w_addr] <= queue_bits_fu_op_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_3_en & queue_bits_wb_id__T_3_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_3_addr] <= queue_bits_wb_id__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_4_en & queue_bits_wb_id__T_4_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_4_addr] <= queue_bits_wb_id__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_5_en & queue_bits_wb_id__T_5_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_5_addr] <= queue_bits_wb_id__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_6_en & queue_bits_wb_id__T_6_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_6_addr] <= queue_bits_wb_id__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_7_en & queue_bits_wb_id__T_7_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_7_addr] <= queue_bits_wb_id__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_8_en & queue_bits_wb_id__T_8_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_8_addr] <= queue_bits_wb_id__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_9_en & queue_bits_wb_id__T_9_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_9_addr] <= queue_bits_wb_id__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_10_en & queue_bits_wb_id__T_10_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_10_addr] <= queue_bits_wb_id__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_11_en & queue_bits_wb_id__T_11_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_11_addr] <= queue_bits_wb_id__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_12_en & queue_bits_wb_id__T_12_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_12_addr] <= queue_bits_wb_id__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_13_en & queue_bits_wb_id__T_13_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_13_addr] <= queue_bits_wb_id__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_14_en & queue_bits_wb_id__T_14_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_14_addr] <= queue_bits_wb_id__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_15_en & queue_bits_wb_id__T_15_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_15_addr] <= queue_bits_wb_id__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_16_en & queue_bits_wb_id__T_16_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_16_addr] <= queue_bits_wb_id__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_17_en & queue_bits_wb_id__T_17_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_17_addr] <= queue_bits_wb_id__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_18_en & queue_bits_wb_id__T_18_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_18_addr] <= queue_bits_wb_id__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_19_en & queue_bits_wb_id__T_19_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_19_addr] <= queue_bits_wb_id__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_20_en & queue_bits_wb_id__T_20_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_20_addr] <= queue_bits_wb_id__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_21_en & queue_bits_wb_id__T_21_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_21_addr] <= queue_bits_wb_id__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_22_en & queue_bits_wb_id__T_22_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_22_addr] <= queue_bits_wb_id__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_23_en & queue_bits_wb_id__T_23_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_23_addr] <= queue_bits_wb_id__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_24_en & queue_bits_wb_id__T_24_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_24_addr] <= queue_bits_wb_id__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_25_en & queue_bits_wb_id__T_25_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_25_addr] <= queue_bits_wb_id__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_26_en & queue_bits_wb_id__T_26_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_26_addr] <= queue_bits_wb_id__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_27_en & queue_bits_wb_id__T_27_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_27_addr] <= queue_bits_wb_id__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_28_en & queue_bits_wb_id__T_28_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_28_addr] <= queue_bits_wb_id__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_29_en & queue_bits_wb_id__T_29_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_29_addr] <= queue_bits_wb_id__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_30_en & queue_bits_wb_id__T_30_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_30_addr] <= queue_bits_wb_id__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_31_en & queue_bits_wb_id__T_31_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_31_addr] <= queue_bits_wb_id__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_32_en & queue_bits_wb_id__T_32_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_32_addr] <= queue_bits_wb_id__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_33_en & queue_bits_wb_id__T_33_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_33_addr] <= queue_bits_wb_id__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_34_en & queue_bits_wb_id__T_34_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_34_addr] <= queue_bits_wb_id__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_35_en & queue_bits_wb_id__T_35_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_35_addr] <= queue_bits_wb_id__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_36_en & queue_bits_wb_id__T_36_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_36_addr] <= queue_bits_wb_id__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_37_en & queue_bits_wb_id__T_37_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_37_addr] <= queue_bits_wb_id__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_38_en & queue_bits_wb_id__T_38_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_38_addr] <= queue_bits_wb_id__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_39_en & queue_bits_wb_id__T_39_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_39_addr] <= queue_bits_wb_id__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_40_en & queue_bits_wb_id__T_40_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_40_addr] <= queue_bits_wb_id__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_41_en & queue_bits_wb_id__T_41_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_41_addr] <= queue_bits_wb_id__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_42_en & queue_bits_wb_id__T_42_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_42_addr] <= queue_bits_wb_id__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_43_en & queue_bits_wb_id__T_43_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_43_addr] <= queue_bits_wb_id__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_44_en & queue_bits_wb_id__T_44_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_44_addr] <= queue_bits_wb_id__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_45_en & queue_bits_wb_id__T_45_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_45_addr] <= queue_bits_wb_id__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_46_en & queue_bits_wb_id__T_46_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_46_addr] <= queue_bits_wb_id__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_47_en & queue_bits_wb_id__T_47_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_47_addr] <= queue_bits_wb_id__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_48_en & queue_bits_wb_id__T_48_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_48_addr] <= queue_bits_wb_id__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_49_en & queue_bits_wb_id__T_49_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_49_addr] <= queue_bits_wb_id__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_50_en & queue_bits_wb_id__T_50_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_50_addr] <= queue_bits_wb_id__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_51_en & queue_bits_wb_id__T_51_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_51_addr] <= queue_bits_wb_id__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_52_en & queue_bits_wb_id__T_52_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_52_addr] <= queue_bits_wb_id__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_53_en & queue_bits_wb_id__T_53_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_53_addr] <= queue_bits_wb_id__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_54_en & queue_bits_wb_id__T_54_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_54_addr] <= queue_bits_wb_id__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_55_en & queue_bits_wb_id__T_55_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_55_addr] <= queue_bits_wb_id__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_56_en & queue_bits_wb_id__T_56_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_56_addr] <= queue_bits_wb_id__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_57_en & queue_bits_wb_id__T_57_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_57_addr] <= queue_bits_wb_id__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_58_en & queue_bits_wb_id__T_58_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_58_addr] <= queue_bits_wb_id__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_59_en & queue_bits_wb_id__T_59_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_59_addr] <= queue_bits_wb_id__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_60_en & queue_bits_wb_id__T_60_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_60_addr] <= queue_bits_wb_id__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_61_en & queue_bits_wb_id__T_61_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_61_addr] <= queue_bits_wb_id__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_62_en & queue_bits_wb_id__T_62_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_62_addr] <= queue_bits_wb_id__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_63_en & queue_bits_wb_id__T_63_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_63_addr] <= queue_bits_wb_id__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_64_en & queue_bits_wb_id__T_64_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_64_addr] <= queue_bits_wb_id__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_65_en & queue_bits_wb_id__T_65_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_65_addr] <= queue_bits_wb_id__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_66_en & queue_bits_wb_id__T_66_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_66_addr] <= queue_bits_wb_id__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_67_en & queue_bits_wb_id__T_67_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_67_addr] <= queue_bits_wb_id__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_68_en & queue_bits_wb_id__T_68_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_68_addr] <= queue_bits_wb_id__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_70_en & queue_bits_wb_id__T_70_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_70_addr] <= queue_bits_wb_id__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_71_en & queue_bits_wb_id__T_71_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_71_addr] <= queue_bits_wb_id__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_72_en & queue_bits_wb_id__T_72_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_72_addr] <= queue_bits_wb_id__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_73_en & queue_bits_wb_id__T_73_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_73_addr] <= queue_bits_wb_id__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_74_en & queue_bits_wb_id__T_74_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_74_addr] <= queue_bits_wb_id__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_75_en & queue_bits_wb_id__T_75_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_75_addr] <= queue_bits_wb_id__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_76_en & queue_bits_wb_id__T_76_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_76_addr] <= queue_bits_wb_id__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_77_en & queue_bits_wb_id__T_77_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_77_addr] <= queue_bits_wb_id__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_78_en & queue_bits_wb_id__T_78_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_78_addr] <= queue_bits_wb_id__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_79_en & queue_bits_wb_id__T_79_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_79_addr] <= queue_bits_wb_id__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_80_en & queue_bits_wb_id__T_80_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_80_addr] <= queue_bits_wb_id__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_81_en & queue_bits_wb_id__T_81_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_81_addr] <= queue_bits_wb_id__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_82_en & queue_bits_wb_id__T_82_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_82_addr] <= queue_bits_wb_id__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_83_en & queue_bits_wb_id__T_83_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_83_addr] <= queue_bits_wb_id__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_84_en & queue_bits_wb_id__T_84_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_84_addr] <= queue_bits_wb_id__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_85_en & queue_bits_wb_id__T_85_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_85_addr] <= queue_bits_wb_id__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_86_en & queue_bits_wb_id__T_86_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_86_addr] <= queue_bits_wb_id__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_87_en & queue_bits_wb_id__T_87_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_87_addr] <= queue_bits_wb_id__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_88_en & queue_bits_wb_id__T_88_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_88_addr] <= queue_bits_wb_id__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_89_en & queue_bits_wb_id__T_89_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_89_addr] <= queue_bits_wb_id__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_90_en & queue_bits_wb_id__T_90_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_90_addr] <= queue_bits_wb_id__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_91_en & queue_bits_wb_id__T_91_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_91_addr] <= queue_bits_wb_id__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_92_en & queue_bits_wb_id__T_92_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_92_addr] <= queue_bits_wb_id__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_93_en & queue_bits_wb_id__T_93_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_93_addr] <= queue_bits_wb_id__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_94_en & queue_bits_wb_id__T_94_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_94_addr] <= queue_bits_wb_id__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_95_en & queue_bits_wb_id__T_95_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_95_addr] <= queue_bits_wb_id__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_96_en & queue_bits_wb_id__T_96_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_96_addr] <= queue_bits_wb_id__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_97_en & queue_bits_wb_id__T_97_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_97_addr] <= queue_bits_wb_id__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_98_en & queue_bits_wb_id__T_98_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_98_addr] <= queue_bits_wb_id__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_99_en & queue_bits_wb_id__T_99_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_99_addr] <= queue_bits_wb_id__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_100_en & queue_bits_wb_id__T_100_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_100_addr] <= queue_bits_wb_id__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_101_en & queue_bits_wb_id__T_101_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_101_addr] <= queue_bits_wb_id__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_102_en & queue_bits_wb_id__T_102_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_102_addr] <= queue_bits_wb_id__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_103_en & queue_bits_wb_id__T_103_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_103_addr] <= queue_bits_wb_id__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_104_en & queue_bits_wb_id__T_104_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_104_addr] <= queue_bits_wb_id__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_105_en & queue_bits_wb_id__T_105_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_105_addr] <= queue_bits_wb_id__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_106_en & queue_bits_wb_id__T_106_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_106_addr] <= queue_bits_wb_id__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_107_en & queue_bits_wb_id__T_107_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_107_addr] <= queue_bits_wb_id__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_108_en & queue_bits_wb_id__T_108_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_108_addr] <= queue_bits_wb_id__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_109_en & queue_bits_wb_id__T_109_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_109_addr] <= queue_bits_wb_id__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_110_en & queue_bits_wb_id__T_110_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_110_addr] <= queue_bits_wb_id__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_111_en & queue_bits_wb_id__T_111_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_111_addr] <= queue_bits_wb_id__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_112_en & queue_bits_wb_id__T_112_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_112_addr] <= queue_bits_wb_id__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_113_en & queue_bits_wb_id__T_113_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_113_addr] <= queue_bits_wb_id__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_114_en & queue_bits_wb_id__T_114_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_114_addr] <= queue_bits_wb_id__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_115_en & queue_bits_wb_id__T_115_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_115_addr] <= queue_bits_wb_id__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_116_en & queue_bits_wb_id__T_116_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_116_addr] <= queue_bits_wb_id__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_117_en & queue_bits_wb_id__T_117_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_117_addr] <= queue_bits_wb_id__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_118_en & queue_bits_wb_id__T_118_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_118_addr] <= queue_bits_wb_id__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_119_en & queue_bits_wb_id__T_119_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_119_addr] <= queue_bits_wb_id__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_120_en & queue_bits_wb_id__T_120_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_120_addr] <= queue_bits_wb_id__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_121_en & queue_bits_wb_id__T_121_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_121_addr] <= queue_bits_wb_id__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_122_en & queue_bits_wb_id__T_122_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_122_addr] <= queue_bits_wb_id__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_123_en & queue_bits_wb_id__T_123_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_123_addr] <= queue_bits_wb_id__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_124_en & queue_bits_wb_id__T_124_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_124_addr] <= queue_bits_wb_id__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_125_en & queue_bits_wb_id__T_125_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_125_addr] <= queue_bits_wb_id__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_126_en & queue_bits_wb_id__T_126_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_126_addr] <= queue_bits_wb_id__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_127_en & queue_bits_wb_id__T_127_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_127_addr] <= queue_bits_wb_id__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_128_en & queue_bits_wb_id__T_128_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_128_addr] <= queue_bits_wb_id__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_129_en & queue_bits_wb_id__T_129_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_129_addr] <= queue_bits_wb_id__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_130_en & queue_bits_wb_id__T_130_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_130_addr] <= queue_bits_wb_id__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_131_en & queue_bits_wb_id__T_131_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_131_addr] <= queue_bits_wb_id__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_132_en & queue_bits_wb_id__T_132_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_132_addr] <= queue_bits_wb_id__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id__T_133_en & queue_bits_wb_id__T_133_mask) begin
      queue_bits_wb_id[queue_bits_wb_id__T_133_addr] <= queue_bits_wb_id__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_id_q_head_w_en & queue_bits_wb_id_q_head_w_mask) begin
      queue_bits_wb_id[queue_bits_wb_id_q_head_w_addr] <= queue_bits_wb_id_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_3_en & queue_bits_wb_pc__T_3_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_3_addr] <= queue_bits_wb_pc__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_4_en & queue_bits_wb_pc__T_4_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_4_addr] <= queue_bits_wb_pc__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_5_en & queue_bits_wb_pc__T_5_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_5_addr] <= queue_bits_wb_pc__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_6_en & queue_bits_wb_pc__T_6_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_6_addr] <= queue_bits_wb_pc__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_7_en & queue_bits_wb_pc__T_7_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_7_addr] <= queue_bits_wb_pc__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_8_en & queue_bits_wb_pc__T_8_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_8_addr] <= queue_bits_wb_pc__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_9_en & queue_bits_wb_pc__T_9_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_9_addr] <= queue_bits_wb_pc__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_10_en & queue_bits_wb_pc__T_10_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_10_addr] <= queue_bits_wb_pc__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_11_en & queue_bits_wb_pc__T_11_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_11_addr] <= queue_bits_wb_pc__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_12_en & queue_bits_wb_pc__T_12_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_12_addr] <= queue_bits_wb_pc__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_13_en & queue_bits_wb_pc__T_13_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_13_addr] <= queue_bits_wb_pc__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_14_en & queue_bits_wb_pc__T_14_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_14_addr] <= queue_bits_wb_pc__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_15_en & queue_bits_wb_pc__T_15_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_15_addr] <= queue_bits_wb_pc__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_16_en & queue_bits_wb_pc__T_16_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_16_addr] <= queue_bits_wb_pc__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_17_en & queue_bits_wb_pc__T_17_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_17_addr] <= queue_bits_wb_pc__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_18_en & queue_bits_wb_pc__T_18_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_18_addr] <= queue_bits_wb_pc__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_19_en & queue_bits_wb_pc__T_19_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_19_addr] <= queue_bits_wb_pc__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_20_en & queue_bits_wb_pc__T_20_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_20_addr] <= queue_bits_wb_pc__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_21_en & queue_bits_wb_pc__T_21_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_21_addr] <= queue_bits_wb_pc__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_22_en & queue_bits_wb_pc__T_22_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_22_addr] <= queue_bits_wb_pc__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_23_en & queue_bits_wb_pc__T_23_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_23_addr] <= queue_bits_wb_pc__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_24_en & queue_bits_wb_pc__T_24_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_24_addr] <= queue_bits_wb_pc__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_25_en & queue_bits_wb_pc__T_25_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_25_addr] <= queue_bits_wb_pc__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_26_en & queue_bits_wb_pc__T_26_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_26_addr] <= queue_bits_wb_pc__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_27_en & queue_bits_wb_pc__T_27_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_27_addr] <= queue_bits_wb_pc__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_28_en & queue_bits_wb_pc__T_28_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_28_addr] <= queue_bits_wb_pc__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_29_en & queue_bits_wb_pc__T_29_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_29_addr] <= queue_bits_wb_pc__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_30_en & queue_bits_wb_pc__T_30_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_30_addr] <= queue_bits_wb_pc__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_31_en & queue_bits_wb_pc__T_31_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_31_addr] <= queue_bits_wb_pc__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_32_en & queue_bits_wb_pc__T_32_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_32_addr] <= queue_bits_wb_pc__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_33_en & queue_bits_wb_pc__T_33_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_33_addr] <= queue_bits_wb_pc__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_34_en & queue_bits_wb_pc__T_34_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_34_addr] <= queue_bits_wb_pc__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_35_en & queue_bits_wb_pc__T_35_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_35_addr] <= queue_bits_wb_pc__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_36_en & queue_bits_wb_pc__T_36_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_36_addr] <= queue_bits_wb_pc__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_37_en & queue_bits_wb_pc__T_37_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_37_addr] <= queue_bits_wb_pc__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_38_en & queue_bits_wb_pc__T_38_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_38_addr] <= queue_bits_wb_pc__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_39_en & queue_bits_wb_pc__T_39_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_39_addr] <= queue_bits_wb_pc__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_40_en & queue_bits_wb_pc__T_40_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_40_addr] <= queue_bits_wb_pc__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_41_en & queue_bits_wb_pc__T_41_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_41_addr] <= queue_bits_wb_pc__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_42_en & queue_bits_wb_pc__T_42_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_42_addr] <= queue_bits_wb_pc__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_43_en & queue_bits_wb_pc__T_43_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_43_addr] <= queue_bits_wb_pc__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_44_en & queue_bits_wb_pc__T_44_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_44_addr] <= queue_bits_wb_pc__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_45_en & queue_bits_wb_pc__T_45_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_45_addr] <= queue_bits_wb_pc__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_46_en & queue_bits_wb_pc__T_46_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_46_addr] <= queue_bits_wb_pc__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_47_en & queue_bits_wb_pc__T_47_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_47_addr] <= queue_bits_wb_pc__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_48_en & queue_bits_wb_pc__T_48_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_48_addr] <= queue_bits_wb_pc__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_49_en & queue_bits_wb_pc__T_49_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_49_addr] <= queue_bits_wb_pc__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_50_en & queue_bits_wb_pc__T_50_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_50_addr] <= queue_bits_wb_pc__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_51_en & queue_bits_wb_pc__T_51_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_51_addr] <= queue_bits_wb_pc__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_52_en & queue_bits_wb_pc__T_52_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_52_addr] <= queue_bits_wb_pc__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_53_en & queue_bits_wb_pc__T_53_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_53_addr] <= queue_bits_wb_pc__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_54_en & queue_bits_wb_pc__T_54_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_54_addr] <= queue_bits_wb_pc__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_55_en & queue_bits_wb_pc__T_55_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_55_addr] <= queue_bits_wb_pc__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_56_en & queue_bits_wb_pc__T_56_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_56_addr] <= queue_bits_wb_pc__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_57_en & queue_bits_wb_pc__T_57_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_57_addr] <= queue_bits_wb_pc__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_58_en & queue_bits_wb_pc__T_58_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_58_addr] <= queue_bits_wb_pc__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_59_en & queue_bits_wb_pc__T_59_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_59_addr] <= queue_bits_wb_pc__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_60_en & queue_bits_wb_pc__T_60_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_60_addr] <= queue_bits_wb_pc__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_61_en & queue_bits_wb_pc__T_61_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_61_addr] <= queue_bits_wb_pc__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_62_en & queue_bits_wb_pc__T_62_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_62_addr] <= queue_bits_wb_pc__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_63_en & queue_bits_wb_pc__T_63_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_63_addr] <= queue_bits_wb_pc__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_64_en & queue_bits_wb_pc__T_64_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_64_addr] <= queue_bits_wb_pc__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_65_en & queue_bits_wb_pc__T_65_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_65_addr] <= queue_bits_wb_pc__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_66_en & queue_bits_wb_pc__T_66_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_66_addr] <= queue_bits_wb_pc__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_67_en & queue_bits_wb_pc__T_67_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_67_addr] <= queue_bits_wb_pc__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_68_en & queue_bits_wb_pc__T_68_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_68_addr] <= queue_bits_wb_pc__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_70_en & queue_bits_wb_pc__T_70_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_70_addr] <= queue_bits_wb_pc__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_71_en & queue_bits_wb_pc__T_71_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_71_addr] <= queue_bits_wb_pc__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_72_en & queue_bits_wb_pc__T_72_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_72_addr] <= queue_bits_wb_pc__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_73_en & queue_bits_wb_pc__T_73_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_73_addr] <= queue_bits_wb_pc__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_74_en & queue_bits_wb_pc__T_74_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_74_addr] <= queue_bits_wb_pc__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_75_en & queue_bits_wb_pc__T_75_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_75_addr] <= queue_bits_wb_pc__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_76_en & queue_bits_wb_pc__T_76_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_76_addr] <= queue_bits_wb_pc__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_77_en & queue_bits_wb_pc__T_77_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_77_addr] <= queue_bits_wb_pc__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_78_en & queue_bits_wb_pc__T_78_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_78_addr] <= queue_bits_wb_pc__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_79_en & queue_bits_wb_pc__T_79_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_79_addr] <= queue_bits_wb_pc__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_80_en & queue_bits_wb_pc__T_80_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_80_addr] <= queue_bits_wb_pc__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_81_en & queue_bits_wb_pc__T_81_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_81_addr] <= queue_bits_wb_pc__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_82_en & queue_bits_wb_pc__T_82_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_82_addr] <= queue_bits_wb_pc__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_83_en & queue_bits_wb_pc__T_83_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_83_addr] <= queue_bits_wb_pc__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_84_en & queue_bits_wb_pc__T_84_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_84_addr] <= queue_bits_wb_pc__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_85_en & queue_bits_wb_pc__T_85_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_85_addr] <= queue_bits_wb_pc__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_86_en & queue_bits_wb_pc__T_86_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_86_addr] <= queue_bits_wb_pc__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_87_en & queue_bits_wb_pc__T_87_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_87_addr] <= queue_bits_wb_pc__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_88_en & queue_bits_wb_pc__T_88_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_88_addr] <= queue_bits_wb_pc__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_89_en & queue_bits_wb_pc__T_89_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_89_addr] <= queue_bits_wb_pc__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_90_en & queue_bits_wb_pc__T_90_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_90_addr] <= queue_bits_wb_pc__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_91_en & queue_bits_wb_pc__T_91_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_91_addr] <= queue_bits_wb_pc__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_92_en & queue_bits_wb_pc__T_92_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_92_addr] <= queue_bits_wb_pc__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_93_en & queue_bits_wb_pc__T_93_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_93_addr] <= queue_bits_wb_pc__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_94_en & queue_bits_wb_pc__T_94_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_94_addr] <= queue_bits_wb_pc__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_95_en & queue_bits_wb_pc__T_95_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_95_addr] <= queue_bits_wb_pc__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_96_en & queue_bits_wb_pc__T_96_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_96_addr] <= queue_bits_wb_pc__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_97_en & queue_bits_wb_pc__T_97_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_97_addr] <= queue_bits_wb_pc__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_98_en & queue_bits_wb_pc__T_98_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_98_addr] <= queue_bits_wb_pc__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_99_en & queue_bits_wb_pc__T_99_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_99_addr] <= queue_bits_wb_pc__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_100_en & queue_bits_wb_pc__T_100_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_100_addr] <= queue_bits_wb_pc__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_101_en & queue_bits_wb_pc__T_101_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_101_addr] <= queue_bits_wb_pc__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_102_en & queue_bits_wb_pc__T_102_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_102_addr] <= queue_bits_wb_pc__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_103_en & queue_bits_wb_pc__T_103_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_103_addr] <= queue_bits_wb_pc__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_104_en & queue_bits_wb_pc__T_104_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_104_addr] <= queue_bits_wb_pc__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_105_en & queue_bits_wb_pc__T_105_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_105_addr] <= queue_bits_wb_pc__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_106_en & queue_bits_wb_pc__T_106_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_106_addr] <= queue_bits_wb_pc__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_107_en & queue_bits_wb_pc__T_107_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_107_addr] <= queue_bits_wb_pc__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_108_en & queue_bits_wb_pc__T_108_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_108_addr] <= queue_bits_wb_pc__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_109_en & queue_bits_wb_pc__T_109_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_109_addr] <= queue_bits_wb_pc__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_110_en & queue_bits_wb_pc__T_110_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_110_addr] <= queue_bits_wb_pc__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_111_en & queue_bits_wb_pc__T_111_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_111_addr] <= queue_bits_wb_pc__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_112_en & queue_bits_wb_pc__T_112_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_112_addr] <= queue_bits_wb_pc__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_113_en & queue_bits_wb_pc__T_113_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_113_addr] <= queue_bits_wb_pc__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_114_en & queue_bits_wb_pc__T_114_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_114_addr] <= queue_bits_wb_pc__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_115_en & queue_bits_wb_pc__T_115_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_115_addr] <= queue_bits_wb_pc__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_116_en & queue_bits_wb_pc__T_116_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_116_addr] <= queue_bits_wb_pc__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_117_en & queue_bits_wb_pc__T_117_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_117_addr] <= queue_bits_wb_pc__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_118_en & queue_bits_wb_pc__T_118_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_118_addr] <= queue_bits_wb_pc__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_119_en & queue_bits_wb_pc__T_119_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_119_addr] <= queue_bits_wb_pc__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_120_en & queue_bits_wb_pc__T_120_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_120_addr] <= queue_bits_wb_pc__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_121_en & queue_bits_wb_pc__T_121_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_121_addr] <= queue_bits_wb_pc__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_122_en & queue_bits_wb_pc__T_122_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_122_addr] <= queue_bits_wb_pc__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_123_en & queue_bits_wb_pc__T_123_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_123_addr] <= queue_bits_wb_pc__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_124_en & queue_bits_wb_pc__T_124_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_124_addr] <= queue_bits_wb_pc__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_125_en & queue_bits_wb_pc__T_125_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_125_addr] <= queue_bits_wb_pc__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_126_en & queue_bits_wb_pc__T_126_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_126_addr] <= queue_bits_wb_pc__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_127_en & queue_bits_wb_pc__T_127_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_127_addr] <= queue_bits_wb_pc__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_128_en & queue_bits_wb_pc__T_128_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_128_addr] <= queue_bits_wb_pc__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_129_en & queue_bits_wb_pc__T_129_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_129_addr] <= queue_bits_wb_pc__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_130_en & queue_bits_wb_pc__T_130_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_130_addr] <= queue_bits_wb_pc__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_131_en & queue_bits_wb_pc__T_131_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_131_addr] <= queue_bits_wb_pc__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_132_en & queue_bits_wb_pc__T_132_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_132_addr] <= queue_bits_wb_pc__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc__T_133_en & queue_bits_wb_pc__T_133_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc__T_133_addr] <= queue_bits_wb_pc__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_pc_q_head_w_en & queue_bits_wb_pc_q_head_w_mask) begin
      queue_bits_wb_pc[queue_bits_wb_pc_q_head_w_addr] <= queue_bits_wb_pc_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_3_en & queue_bits_wb_instr_op__T_3_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_3_addr] <= queue_bits_wb_instr_op__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_4_en & queue_bits_wb_instr_op__T_4_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_4_addr] <= queue_bits_wb_instr_op__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_5_en & queue_bits_wb_instr_op__T_5_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_5_addr] <= queue_bits_wb_instr_op__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_6_en & queue_bits_wb_instr_op__T_6_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_6_addr] <= queue_bits_wb_instr_op__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_7_en & queue_bits_wb_instr_op__T_7_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_7_addr] <= queue_bits_wb_instr_op__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_8_en & queue_bits_wb_instr_op__T_8_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_8_addr] <= queue_bits_wb_instr_op__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_9_en & queue_bits_wb_instr_op__T_9_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_9_addr] <= queue_bits_wb_instr_op__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_10_en & queue_bits_wb_instr_op__T_10_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_10_addr] <= queue_bits_wb_instr_op__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_11_en & queue_bits_wb_instr_op__T_11_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_11_addr] <= queue_bits_wb_instr_op__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_12_en & queue_bits_wb_instr_op__T_12_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_12_addr] <= queue_bits_wb_instr_op__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_13_en & queue_bits_wb_instr_op__T_13_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_13_addr] <= queue_bits_wb_instr_op__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_14_en & queue_bits_wb_instr_op__T_14_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_14_addr] <= queue_bits_wb_instr_op__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_15_en & queue_bits_wb_instr_op__T_15_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_15_addr] <= queue_bits_wb_instr_op__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_16_en & queue_bits_wb_instr_op__T_16_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_16_addr] <= queue_bits_wb_instr_op__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_17_en & queue_bits_wb_instr_op__T_17_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_17_addr] <= queue_bits_wb_instr_op__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_18_en & queue_bits_wb_instr_op__T_18_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_18_addr] <= queue_bits_wb_instr_op__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_19_en & queue_bits_wb_instr_op__T_19_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_19_addr] <= queue_bits_wb_instr_op__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_20_en & queue_bits_wb_instr_op__T_20_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_20_addr] <= queue_bits_wb_instr_op__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_21_en & queue_bits_wb_instr_op__T_21_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_21_addr] <= queue_bits_wb_instr_op__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_22_en & queue_bits_wb_instr_op__T_22_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_22_addr] <= queue_bits_wb_instr_op__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_23_en & queue_bits_wb_instr_op__T_23_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_23_addr] <= queue_bits_wb_instr_op__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_24_en & queue_bits_wb_instr_op__T_24_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_24_addr] <= queue_bits_wb_instr_op__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_25_en & queue_bits_wb_instr_op__T_25_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_25_addr] <= queue_bits_wb_instr_op__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_26_en & queue_bits_wb_instr_op__T_26_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_26_addr] <= queue_bits_wb_instr_op__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_27_en & queue_bits_wb_instr_op__T_27_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_27_addr] <= queue_bits_wb_instr_op__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_28_en & queue_bits_wb_instr_op__T_28_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_28_addr] <= queue_bits_wb_instr_op__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_29_en & queue_bits_wb_instr_op__T_29_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_29_addr] <= queue_bits_wb_instr_op__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_30_en & queue_bits_wb_instr_op__T_30_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_30_addr] <= queue_bits_wb_instr_op__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_31_en & queue_bits_wb_instr_op__T_31_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_31_addr] <= queue_bits_wb_instr_op__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_32_en & queue_bits_wb_instr_op__T_32_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_32_addr] <= queue_bits_wb_instr_op__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_33_en & queue_bits_wb_instr_op__T_33_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_33_addr] <= queue_bits_wb_instr_op__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_34_en & queue_bits_wb_instr_op__T_34_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_34_addr] <= queue_bits_wb_instr_op__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_35_en & queue_bits_wb_instr_op__T_35_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_35_addr] <= queue_bits_wb_instr_op__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_36_en & queue_bits_wb_instr_op__T_36_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_36_addr] <= queue_bits_wb_instr_op__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_37_en & queue_bits_wb_instr_op__T_37_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_37_addr] <= queue_bits_wb_instr_op__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_38_en & queue_bits_wb_instr_op__T_38_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_38_addr] <= queue_bits_wb_instr_op__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_39_en & queue_bits_wb_instr_op__T_39_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_39_addr] <= queue_bits_wb_instr_op__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_40_en & queue_bits_wb_instr_op__T_40_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_40_addr] <= queue_bits_wb_instr_op__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_41_en & queue_bits_wb_instr_op__T_41_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_41_addr] <= queue_bits_wb_instr_op__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_42_en & queue_bits_wb_instr_op__T_42_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_42_addr] <= queue_bits_wb_instr_op__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_43_en & queue_bits_wb_instr_op__T_43_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_43_addr] <= queue_bits_wb_instr_op__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_44_en & queue_bits_wb_instr_op__T_44_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_44_addr] <= queue_bits_wb_instr_op__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_45_en & queue_bits_wb_instr_op__T_45_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_45_addr] <= queue_bits_wb_instr_op__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_46_en & queue_bits_wb_instr_op__T_46_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_46_addr] <= queue_bits_wb_instr_op__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_47_en & queue_bits_wb_instr_op__T_47_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_47_addr] <= queue_bits_wb_instr_op__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_48_en & queue_bits_wb_instr_op__T_48_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_48_addr] <= queue_bits_wb_instr_op__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_49_en & queue_bits_wb_instr_op__T_49_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_49_addr] <= queue_bits_wb_instr_op__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_50_en & queue_bits_wb_instr_op__T_50_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_50_addr] <= queue_bits_wb_instr_op__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_51_en & queue_bits_wb_instr_op__T_51_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_51_addr] <= queue_bits_wb_instr_op__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_52_en & queue_bits_wb_instr_op__T_52_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_52_addr] <= queue_bits_wb_instr_op__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_53_en & queue_bits_wb_instr_op__T_53_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_53_addr] <= queue_bits_wb_instr_op__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_54_en & queue_bits_wb_instr_op__T_54_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_54_addr] <= queue_bits_wb_instr_op__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_55_en & queue_bits_wb_instr_op__T_55_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_55_addr] <= queue_bits_wb_instr_op__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_56_en & queue_bits_wb_instr_op__T_56_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_56_addr] <= queue_bits_wb_instr_op__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_57_en & queue_bits_wb_instr_op__T_57_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_57_addr] <= queue_bits_wb_instr_op__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_58_en & queue_bits_wb_instr_op__T_58_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_58_addr] <= queue_bits_wb_instr_op__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_59_en & queue_bits_wb_instr_op__T_59_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_59_addr] <= queue_bits_wb_instr_op__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_60_en & queue_bits_wb_instr_op__T_60_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_60_addr] <= queue_bits_wb_instr_op__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_61_en & queue_bits_wb_instr_op__T_61_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_61_addr] <= queue_bits_wb_instr_op__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_62_en & queue_bits_wb_instr_op__T_62_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_62_addr] <= queue_bits_wb_instr_op__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_63_en & queue_bits_wb_instr_op__T_63_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_63_addr] <= queue_bits_wb_instr_op__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_64_en & queue_bits_wb_instr_op__T_64_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_64_addr] <= queue_bits_wb_instr_op__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_65_en & queue_bits_wb_instr_op__T_65_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_65_addr] <= queue_bits_wb_instr_op__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_66_en & queue_bits_wb_instr_op__T_66_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_66_addr] <= queue_bits_wb_instr_op__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_67_en & queue_bits_wb_instr_op__T_67_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_67_addr] <= queue_bits_wb_instr_op__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_68_en & queue_bits_wb_instr_op__T_68_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_68_addr] <= queue_bits_wb_instr_op__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_70_en & queue_bits_wb_instr_op__T_70_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_70_addr] <= queue_bits_wb_instr_op__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_71_en & queue_bits_wb_instr_op__T_71_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_71_addr] <= queue_bits_wb_instr_op__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_72_en & queue_bits_wb_instr_op__T_72_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_72_addr] <= queue_bits_wb_instr_op__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_73_en & queue_bits_wb_instr_op__T_73_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_73_addr] <= queue_bits_wb_instr_op__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_74_en & queue_bits_wb_instr_op__T_74_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_74_addr] <= queue_bits_wb_instr_op__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_75_en & queue_bits_wb_instr_op__T_75_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_75_addr] <= queue_bits_wb_instr_op__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_76_en & queue_bits_wb_instr_op__T_76_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_76_addr] <= queue_bits_wb_instr_op__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_77_en & queue_bits_wb_instr_op__T_77_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_77_addr] <= queue_bits_wb_instr_op__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_78_en & queue_bits_wb_instr_op__T_78_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_78_addr] <= queue_bits_wb_instr_op__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_79_en & queue_bits_wb_instr_op__T_79_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_79_addr] <= queue_bits_wb_instr_op__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_80_en & queue_bits_wb_instr_op__T_80_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_80_addr] <= queue_bits_wb_instr_op__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_81_en & queue_bits_wb_instr_op__T_81_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_81_addr] <= queue_bits_wb_instr_op__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_82_en & queue_bits_wb_instr_op__T_82_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_82_addr] <= queue_bits_wb_instr_op__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_83_en & queue_bits_wb_instr_op__T_83_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_83_addr] <= queue_bits_wb_instr_op__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_84_en & queue_bits_wb_instr_op__T_84_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_84_addr] <= queue_bits_wb_instr_op__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_85_en & queue_bits_wb_instr_op__T_85_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_85_addr] <= queue_bits_wb_instr_op__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_86_en & queue_bits_wb_instr_op__T_86_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_86_addr] <= queue_bits_wb_instr_op__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_87_en & queue_bits_wb_instr_op__T_87_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_87_addr] <= queue_bits_wb_instr_op__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_88_en & queue_bits_wb_instr_op__T_88_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_88_addr] <= queue_bits_wb_instr_op__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_89_en & queue_bits_wb_instr_op__T_89_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_89_addr] <= queue_bits_wb_instr_op__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_90_en & queue_bits_wb_instr_op__T_90_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_90_addr] <= queue_bits_wb_instr_op__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_91_en & queue_bits_wb_instr_op__T_91_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_91_addr] <= queue_bits_wb_instr_op__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_92_en & queue_bits_wb_instr_op__T_92_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_92_addr] <= queue_bits_wb_instr_op__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_93_en & queue_bits_wb_instr_op__T_93_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_93_addr] <= queue_bits_wb_instr_op__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_94_en & queue_bits_wb_instr_op__T_94_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_94_addr] <= queue_bits_wb_instr_op__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_95_en & queue_bits_wb_instr_op__T_95_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_95_addr] <= queue_bits_wb_instr_op__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_96_en & queue_bits_wb_instr_op__T_96_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_96_addr] <= queue_bits_wb_instr_op__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_97_en & queue_bits_wb_instr_op__T_97_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_97_addr] <= queue_bits_wb_instr_op__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_98_en & queue_bits_wb_instr_op__T_98_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_98_addr] <= queue_bits_wb_instr_op__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_99_en & queue_bits_wb_instr_op__T_99_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_99_addr] <= queue_bits_wb_instr_op__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_100_en & queue_bits_wb_instr_op__T_100_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_100_addr] <= queue_bits_wb_instr_op__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_101_en & queue_bits_wb_instr_op__T_101_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_101_addr] <= queue_bits_wb_instr_op__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_102_en & queue_bits_wb_instr_op__T_102_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_102_addr] <= queue_bits_wb_instr_op__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_103_en & queue_bits_wb_instr_op__T_103_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_103_addr] <= queue_bits_wb_instr_op__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_104_en & queue_bits_wb_instr_op__T_104_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_104_addr] <= queue_bits_wb_instr_op__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_105_en & queue_bits_wb_instr_op__T_105_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_105_addr] <= queue_bits_wb_instr_op__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_106_en & queue_bits_wb_instr_op__T_106_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_106_addr] <= queue_bits_wb_instr_op__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_107_en & queue_bits_wb_instr_op__T_107_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_107_addr] <= queue_bits_wb_instr_op__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_108_en & queue_bits_wb_instr_op__T_108_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_108_addr] <= queue_bits_wb_instr_op__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_109_en & queue_bits_wb_instr_op__T_109_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_109_addr] <= queue_bits_wb_instr_op__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_110_en & queue_bits_wb_instr_op__T_110_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_110_addr] <= queue_bits_wb_instr_op__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_111_en & queue_bits_wb_instr_op__T_111_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_111_addr] <= queue_bits_wb_instr_op__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_112_en & queue_bits_wb_instr_op__T_112_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_112_addr] <= queue_bits_wb_instr_op__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_113_en & queue_bits_wb_instr_op__T_113_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_113_addr] <= queue_bits_wb_instr_op__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_114_en & queue_bits_wb_instr_op__T_114_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_114_addr] <= queue_bits_wb_instr_op__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_115_en & queue_bits_wb_instr_op__T_115_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_115_addr] <= queue_bits_wb_instr_op__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_116_en & queue_bits_wb_instr_op__T_116_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_116_addr] <= queue_bits_wb_instr_op__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_117_en & queue_bits_wb_instr_op__T_117_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_117_addr] <= queue_bits_wb_instr_op__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_118_en & queue_bits_wb_instr_op__T_118_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_118_addr] <= queue_bits_wb_instr_op__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_119_en & queue_bits_wb_instr_op__T_119_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_119_addr] <= queue_bits_wb_instr_op__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_120_en & queue_bits_wb_instr_op__T_120_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_120_addr] <= queue_bits_wb_instr_op__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_121_en & queue_bits_wb_instr_op__T_121_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_121_addr] <= queue_bits_wb_instr_op__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_122_en & queue_bits_wb_instr_op__T_122_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_122_addr] <= queue_bits_wb_instr_op__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_123_en & queue_bits_wb_instr_op__T_123_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_123_addr] <= queue_bits_wb_instr_op__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_124_en & queue_bits_wb_instr_op__T_124_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_124_addr] <= queue_bits_wb_instr_op__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_125_en & queue_bits_wb_instr_op__T_125_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_125_addr] <= queue_bits_wb_instr_op__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_126_en & queue_bits_wb_instr_op__T_126_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_126_addr] <= queue_bits_wb_instr_op__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_127_en & queue_bits_wb_instr_op__T_127_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_127_addr] <= queue_bits_wb_instr_op__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_128_en & queue_bits_wb_instr_op__T_128_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_128_addr] <= queue_bits_wb_instr_op__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_129_en & queue_bits_wb_instr_op__T_129_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_129_addr] <= queue_bits_wb_instr_op__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_130_en & queue_bits_wb_instr_op__T_130_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_130_addr] <= queue_bits_wb_instr_op__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_131_en & queue_bits_wb_instr_op__T_131_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_131_addr] <= queue_bits_wb_instr_op__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_132_en & queue_bits_wb_instr_op__T_132_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_132_addr] <= queue_bits_wb_instr_op__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op__T_133_en & queue_bits_wb_instr_op__T_133_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op__T_133_addr] <= queue_bits_wb_instr_op__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_op_q_head_w_en & queue_bits_wb_instr_op_q_head_w_mask) begin
      queue_bits_wb_instr_op[queue_bits_wb_instr_op_q_head_w_addr] <= queue_bits_wb_instr_op_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_3_en & queue_bits_wb_instr_rs_idx__T_3_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_3_addr] <= queue_bits_wb_instr_rs_idx__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_4_en & queue_bits_wb_instr_rs_idx__T_4_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_4_addr] <= queue_bits_wb_instr_rs_idx__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_5_en & queue_bits_wb_instr_rs_idx__T_5_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_5_addr] <= queue_bits_wb_instr_rs_idx__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_6_en & queue_bits_wb_instr_rs_idx__T_6_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_6_addr] <= queue_bits_wb_instr_rs_idx__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_7_en & queue_bits_wb_instr_rs_idx__T_7_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_7_addr] <= queue_bits_wb_instr_rs_idx__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_8_en & queue_bits_wb_instr_rs_idx__T_8_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_8_addr] <= queue_bits_wb_instr_rs_idx__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_9_en & queue_bits_wb_instr_rs_idx__T_9_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_9_addr] <= queue_bits_wb_instr_rs_idx__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_10_en & queue_bits_wb_instr_rs_idx__T_10_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_10_addr] <= queue_bits_wb_instr_rs_idx__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_11_en & queue_bits_wb_instr_rs_idx__T_11_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_11_addr] <= queue_bits_wb_instr_rs_idx__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_12_en & queue_bits_wb_instr_rs_idx__T_12_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_12_addr] <= queue_bits_wb_instr_rs_idx__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_13_en & queue_bits_wb_instr_rs_idx__T_13_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_13_addr] <= queue_bits_wb_instr_rs_idx__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_14_en & queue_bits_wb_instr_rs_idx__T_14_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_14_addr] <= queue_bits_wb_instr_rs_idx__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_15_en & queue_bits_wb_instr_rs_idx__T_15_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_15_addr] <= queue_bits_wb_instr_rs_idx__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_16_en & queue_bits_wb_instr_rs_idx__T_16_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_16_addr] <= queue_bits_wb_instr_rs_idx__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_17_en & queue_bits_wb_instr_rs_idx__T_17_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_17_addr] <= queue_bits_wb_instr_rs_idx__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_18_en & queue_bits_wb_instr_rs_idx__T_18_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_18_addr] <= queue_bits_wb_instr_rs_idx__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_19_en & queue_bits_wb_instr_rs_idx__T_19_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_19_addr] <= queue_bits_wb_instr_rs_idx__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_20_en & queue_bits_wb_instr_rs_idx__T_20_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_20_addr] <= queue_bits_wb_instr_rs_idx__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_21_en & queue_bits_wb_instr_rs_idx__T_21_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_21_addr] <= queue_bits_wb_instr_rs_idx__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_22_en & queue_bits_wb_instr_rs_idx__T_22_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_22_addr] <= queue_bits_wb_instr_rs_idx__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_23_en & queue_bits_wb_instr_rs_idx__T_23_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_23_addr] <= queue_bits_wb_instr_rs_idx__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_24_en & queue_bits_wb_instr_rs_idx__T_24_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_24_addr] <= queue_bits_wb_instr_rs_idx__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_25_en & queue_bits_wb_instr_rs_idx__T_25_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_25_addr] <= queue_bits_wb_instr_rs_idx__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_26_en & queue_bits_wb_instr_rs_idx__T_26_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_26_addr] <= queue_bits_wb_instr_rs_idx__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_27_en & queue_bits_wb_instr_rs_idx__T_27_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_27_addr] <= queue_bits_wb_instr_rs_idx__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_28_en & queue_bits_wb_instr_rs_idx__T_28_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_28_addr] <= queue_bits_wb_instr_rs_idx__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_29_en & queue_bits_wb_instr_rs_idx__T_29_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_29_addr] <= queue_bits_wb_instr_rs_idx__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_30_en & queue_bits_wb_instr_rs_idx__T_30_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_30_addr] <= queue_bits_wb_instr_rs_idx__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_31_en & queue_bits_wb_instr_rs_idx__T_31_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_31_addr] <= queue_bits_wb_instr_rs_idx__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_32_en & queue_bits_wb_instr_rs_idx__T_32_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_32_addr] <= queue_bits_wb_instr_rs_idx__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_33_en & queue_bits_wb_instr_rs_idx__T_33_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_33_addr] <= queue_bits_wb_instr_rs_idx__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_34_en & queue_bits_wb_instr_rs_idx__T_34_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_34_addr] <= queue_bits_wb_instr_rs_idx__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_35_en & queue_bits_wb_instr_rs_idx__T_35_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_35_addr] <= queue_bits_wb_instr_rs_idx__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_36_en & queue_bits_wb_instr_rs_idx__T_36_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_36_addr] <= queue_bits_wb_instr_rs_idx__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_37_en & queue_bits_wb_instr_rs_idx__T_37_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_37_addr] <= queue_bits_wb_instr_rs_idx__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_38_en & queue_bits_wb_instr_rs_idx__T_38_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_38_addr] <= queue_bits_wb_instr_rs_idx__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_39_en & queue_bits_wb_instr_rs_idx__T_39_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_39_addr] <= queue_bits_wb_instr_rs_idx__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_40_en & queue_bits_wb_instr_rs_idx__T_40_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_40_addr] <= queue_bits_wb_instr_rs_idx__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_41_en & queue_bits_wb_instr_rs_idx__T_41_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_41_addr] <= queue_bits_wb_instr_rs_idx__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_42_en & queue_bits_wb_instr_rs_idx__T_42_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_42_addr] <= queue_bits_wb_instr_rs_idx__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_43_en & queue_bits_wb_instr_rs_idx__T_43_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_43_addr] <= queue_bits_wb_instr_rs_idx__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_44_en & queue_bits_wb_instr_rs_idx__T_44_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_44_addr] <= queue_bits_wb_instr_rs_idx__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_45_en & queue_bits_wb_instr_rs_idx__T_45_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_45_addr] <= queue_bits_wb_instr_rs_idx__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_46_en & queue_bits_wb_instr_rs_idx__T_46_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_46_addr] <= queue_bits_wb_instr_rs_idx__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_47_en & queue_bits_wb_instr_rs_idx__T_47_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_47_addr] <= queue_bits_wb_instr_rs_idx__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_48_en & queue_bits_wb_instr_rs_idx__T_48_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_48_addr] <= queue_bits_wb_instr_rs_idx__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_49_en & queue_bits_wb_instr_rs_idx__T_49_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_49_addr] <= queue_bits_wb_instr_rs_idx__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_50_en & queue_bits_wb_instr_rs_idx__T_50_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_50_addr] <= queue_bits_wb_instr_rs_idx__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_51_en & queue_bits_wb_instr_rs_idx__T_51_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_51_addr] <= queue_bits_wb_instr_rs_idx__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_52_en & queue_bits_wb_instr_rs_idx__T_52_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_52_addr] <= queue_bits_wb_instr_rs_idx__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_53_en & queue_bits_wb_instr_rs_idx__T_53_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_53_addr] <= queue_bits_wb_instr_rs_idx__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_54_en & queue_bits_wb_instr_rs_idx__T_54_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_54_addr] <= queue_bits_wb_instr_rs_idx__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_55_en & queue_bits_wb_instr_rs_idx__T_55_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_55_addr] <= queue_bits_wb_instr_rs_idx__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_56_en & queue_bits_wb_instr_rs_idx__T_56_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_56_addr] <= queue_bits_wb_instr_rs_idx__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_57_en & queue_bits_wb_instr_rs_idx__T_57_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_57_addr] <= queue_bits_wb_instr_rs_idx__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_58_en & queue_bits_wb_instr_rs_idx__T_58_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_58_addr] <= queue_bits_wb_instr_rs_idx__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_59_en & queue_bits_wb_instr_rs_idx__T_59_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_59_addr] <= queue_bits_wb_instr_rs_idx__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_60_en & queue_bits_wb_instr_rs_idx__T_60_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_60_addr] <= queue_bits_wb_instr_rs_idx__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_61_en & queue_bits_wb_instr_rs_idx__T_61_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_61_addr] <= queue_bits_wb_instr_rs_idx__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_62_en & queue_bits_wb_instr_rs_idx__T_62_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_62_addr] <= queue_bits_wb_instr_rs_idx__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_63_en & queue_bits_wb_instr_rs_idx__T_63_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_63_addr] <= queue_bits_wb_instr_rs_idx__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_64_en & queue_bits_wb_instr_rs_idx__T_64_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_64_addr] <= queue_bits_wb_instr_rs_idx__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_65_en & queue_bits_wb_instr_rs_idx__T_65_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_65_addr] <= queue_bits_wb_instr_rs_idx__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_66_en & queue_bits_wb_instr_rs_idx__T_66_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_66_addr] <= queue_bits_wb_instr_rs_idx__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_67_en & queue_bits_wb_instr_rs_idx__T_67_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_67_addr] <= queue_bits_wb_instr_rs_idx__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_68_en & queue_bits_wb_instr_rs_idx__T_68_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_68_addr] <= queue_bits_wb_instr_rs_idx__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_70_en & queue_bits_wb_instr_rs_idx__T_70_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_70_addr] <= queue_bits_wb_instr_rs_idx__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_71_en & queue_bits_wb_instr_rs_idx__T_71_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_71_addr] <= queue_bits_wb_instr_rs_idx__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_72_en & queue_bits_wb_instr_rs_idx__T_72_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_72_addr] <= queue_bits_wb_instr_rs_idx__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_73_en & queue_bits_wb_instr_rs_idx__T_73_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_73_addr] <= queue_bits_wb_instr_rs_idx__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_74_en & queue_bits_wb_instr_rs_idx__T_74_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_74_addr] <= queue_bits_wb_instr_rs_idx__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_75_en & queue_bits_wb_instr_rs_idx__T_75_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_75_addr] <= queue_bits_wb_instr_rs_idx__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_76_en & queue_bits_wb_instr_rs_idx__T_76_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_76_addr] <= queue_bits_wb_instr_rs_idx__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_77_en & queue_bits_wb_instr_rs_idx__T_77_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_77_addr] <= queue_bits_wb_instr_rs_idx__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_78_en & queue_bits_wb_instr_rs_idx__T_78_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_78_addr] <= queue_bits_wb_instr_rs_idx__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_79_en & queue_bits_wb_instr_rs_idx__T_79_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_79_addr] <= queue_bits_wb_instr_rs_idx__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_80_en & queue_bits_wb_instr_rs_idx__T_80_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_80_addr] <= queue_bits_wb_instr_rs_idx__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_81_en & queue_bits_wb_instr_rs_idx__T_81_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_81_addr] <= queue_bits_wb_instr_rs_idx__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_82_en & queue_bits_wb_instr_rs_idx__T_82_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_82_addr] <= queue_bits_wb_instr_rs_idx__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_83_en & queue_bits_wb_instr_rs_idx__T_83_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_83_addr] <= queue_bits_wb_instr_rs_idx__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_84_en & queue_bits_wb_instr_rs_idx__T_84_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_84_addr] <= queue_bits_wb_instr_rs_idx__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_85_en & queue_bits_wb_instr_rs_idx__T_85_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_85_addr] <= queue_bits_wb_instr_rs_idx__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_86_en & queue_bits_wb_instr_rs_idx__T_86_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_86_addr] <= queue_bits_wb_instr_rs_idx__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_87_en & queue_bits_wb_instr_rs_idx__T_87_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_87_addr] <= queue_bits_wb_instr_rs_idx__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_88_en & queue_bits_wb_instr_rs_idx__T_88_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_88_addr] <= queue_bits_wb_instr_rs_idx__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_89_en & queue_bits_wb_instr_rs_idx__T_89_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_89_addr] <= queue_bits_wb_instr_rs_idx__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_90_en & queue_bits_wb_instr_rs_idx__T_90_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_90_addr] <= queue_bits_wb_instr_rs_idx__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_91_en & queue_bits_wb_instr_rs_idx__T_91_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_91_addr] <= queue_bits_wb_instr_rs_idx__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_92_en & queue_bits_wb_instr_rs_idx__T_92_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_92_addr] <= queue_bits_wb_instr_rs_idx__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_93_en & queue_bits_wb_instr_rs_idx__T_93_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_93_addr] <= queue_bits_wb_instr_rs_idx__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_94_en & queue_bits_wb_instr_rs_idx__T_94_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_94_addr] <= queue_bits_wb_instr_rs_idx__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_95_en & queue_bits_wb_instr_rs_idx__T_95_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_95_addr] <= queue_bits_wb_instr_rs_idx__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_96_en & queue_bits_wb_instr_rs_idx__T_96_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_96_addr] <= queue_bits_wb_instr_rs_idx__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_97_en & queue_bits_wb_instr_rs_idx__T_97_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_97_addr] <= queue_bits_wb_instr_rs_idx__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_98_en & queue_bits_wb_instr_rs_idx__T_98_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_98_addr] <= queue_bits_wb_instr_rs_idx__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_99_en & queue_bits_wb_instr_rs_idx__T_99_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_99_addr] <= queue_bits_wb_instr_rs_idx__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_100_en & queue_bits_wb_instr_rs_idx__T_100_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_100_addr] <= queue_bits_wb_instr_rs_idx__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_101_en & queue_bits_wb_instr_rs_idx__T_101_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_101_addr] <= queue_bits_wb_instr_rs_idx__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_102_en & queue_bits_wb_instr_rs_idx__T_102_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_102_addr] <= queue_bits_wb_instr_rs_idx__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_103_en & queue_bits_wb_instr_rs_idx__T_103_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_103_addr] <= queue_bits_wb_instr_rs_idx__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_104_en & queue_bits_wb_instr_rs_idx__T_104_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_104_addr] <= queue_bits_wb_instr_rs_idx__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_105_en & queue_bits_wb_instr_rs_idx__T_105_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_105_addr] <= queue_bits_wb_instr_rs_idx__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_106_en & queue_bits_wb_instr_rs_idx__T_106_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_106_addr] <= queue_bits_wb_instr_rs_idx__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_107_en & queue_bits_wb_instr_rs_idx__T_107_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_107_addr] <= queue_bits_wb_instr_rs_idx__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_108_en & queue_bits_wb_instr_rs_idx__T_108_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_108_addr] <= queue_bits_wb_instr_rs_idx__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_109_en & queue_bits_wb_instr_rs_idx__T_109_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_109_addr] <= queue_bits_wb_instr_rs_idx__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_110_en & queue_bits_wb_instr_rs_idx__T_110_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_110_addr] <= queue_bits_wb_instr_rs_idx__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_111_en & queue_bits_wb_instr_rs_idx__T_111_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_111_addr] <= queue_bits_wb_instr_rs_idx__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_112_en & queue_bits_wb_instr_rs_idx__T_112_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_112_addr] <= queue_bits_wb_instr_rs_idx__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_113_en & queue_bits_wb_instr_rs_idx__T_113_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_113_addr] <= queue_bits_wb_instr_rs_idx__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_114_en & queue_bits_wb_instr_rs_idx__T_114_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_114_addr] <= queue_bits_wb_instr_rs_idx__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_115_en & queue_bits_wb_instr_rs_idx__T_115_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_115_addr] <= queue_bits_wb_instr_rs_idx__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_116_en & queue_bits_wb_instr_rs_idx__T_116_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_116_addr] <= queue_bits_wb_instr_rs_idx__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_117_en & queue_bits_wb_instr_rs_idx__T_117_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_117_addr] <= queue_bits_wb_instr_rs_idx__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_118_en & queue_bits_wb_instr_rs_idx__T_118_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_118_addr] <= queue_bits_wb_instr_rs_idx__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_119_en & queue_bits_wb_instr_rs_idx__T_119_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_119_addr] <= queue_bits_wb_instr_rs_idx__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_120_en & queue_bits_wb_instr_rs_idx__T_120_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_120_addr] <= queue_bits_wb_instr_rs_idx__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_121_en & queue_bits_wb_instr_rs_idx__T_121_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_121_addr] <= queue_bits_wb_instr_rs_idx__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_122_en & queue_bits_wb_instr_rs_idx__T_122_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_122_addr] <= queue_bits_wb_instr_rs_idx__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_123_en & queue_bits_wb_instr_rs_idx__T_123_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_123_addr] <= queue_bits_wb_instr_rs_idx__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_124_en & queue_bits_wb_instr_rs_idx__T_124_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_124_addr] <= queue_bits_wb_instr_rs_idx__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_125_en & queue_bits_wb_instr_rs_idx__T_125_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_125_addr] <= queue_bits_wb_instr_rs_idx__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_126_en & queue_bits_wb_instr_rs_idx__T_126_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_126_addr] <= queue_bits_wb_instr_rs_idx__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_127_en & queue_bits_wb_instr_rs_idx__T_127_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_127_addr] <= queue_bits_wb_instr_rs_idx__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_128_en & queue_bits_wb_instr_rs_idx__T_128_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_128_addr] <= queue_bits_wb_instr_rs_idx__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_129_en & queue_bits_wb_instr_rs_idx__T_129_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_129_addr] <= queue_bits_wb_instr_rs_idx__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_130_en & queue_bits_wb_instr_rs_idx__T_130_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_130_addr] <= queue_bits_wb_instr_rs_idx__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_131_en & queue_bits_wb_instr_rs_idx__T_131_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_131_addr] <= queue_bits_wb_instr_rs_idx__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_132_en & queue_bits_wb_instr_rs_idx__T_132_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_132_addr] <= queue_bits_wb_instr_rs_idx__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx__T_133_en & queue_bits_wb_instr_rs_idx__T_133_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx__T_133_addr] <= queue_bits_wb_instr_rs_idx__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rs_idx_q_head_w_en & queue_bits_wb_instr_rs_idx_q_head_w_mask) begin
      queue_bits_wb_instr_rs_idx[queue_bits_wb_instr_rs_idx_q_head_w_addr] <= queue_bits_wb_instr_rs_idx_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_3_en & queue_bits_wb_instr_rt_idx__T_3_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_3_addr] <= queue_bits_wb_instr_rt_idx__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_4_en & queue_bits_wb_instr_rt_idx__T_4_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_4_addr] <= queue_bits_wb_instr_rt_idx__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_5_en & queue_bits_wb_instr_rt_idx__T_5_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_5_addr] <= queue_bits_wb_instr_rt_idx__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_6_en & queue_bits_wb_instr_rt_idx__T_6_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_6_addr] <= queue_bits_wb_instr_rt_idx__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_7_en & queue_bits_wb_instr_rt_idx__T_7_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_7_addr] <= queue_bits_wb_instr_rt_idx__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_8_en & queue_bits_wb_instr_rt_idx__T_8_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_8_addr] <= queue_bits_wb_instr_rt_idx__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_9_en & queue_bits_wb_instr_rt_idx__T_9_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_9_addr] <= queue_bits_wb_instr_rt_idx__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_10_en & queue_bits_wb_instr_rt_idx__T_10_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_10_addr] <= queue_bits_wb_instr_rt_idx__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_11_en & queue_bits_wb_instr_rt_idx__T_11_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_11_addr] <= queue_bits_wb_instr_rt_idx__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_12_en & queue_bits_wb_instr_rt_idx__T_12_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_12_addr] <= queue_bits_wb_instr_rt_idx__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_13_en & queue_bits_wb_instr_rt_idx__T_13_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_13_addr] <= queue_bits_wb_instr_rt_idx__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_14_en & queue_bits_wb_instr_rt_idx__T_14_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_14_addr] <= queue_bits_wb_instr_rt_idx__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_15_en & queue_bits_wb_instr_rt_idx__T_15_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_15_addr] <= queue_bits_wb_instr_rt_idx__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_16_en & queue_bits_wb_instr_rt_idx__T_16_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_16_addr] <= queue_bits_wb_instr_rt_idx__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_17_en & queue_bits_wb_instr_rt_idx__T_17_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_17_addr] <= queue_bits_wb_instr_rt_idx__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_18_en & queue_bits_wb_instr_rt_idx__T_18_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_18_addr] <= queue_bits_wb_instr_rt_idx__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_19_en & queue_bits_wb_instr_rt_idx__T_19_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_19_addr] <= queue_bits_wb_instr_rt_idx__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_20_en & queue_bits_wb_instr_rt_idx__T_20_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_20_addr] <= queue_bits_wb_instr_rt_idx__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_21_en & queue_bits_wb_instr_rt_idx__T_21_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_21_addr] <= queue_bits_wb_instr_rt_idx__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_22_en & queue_bits_wb_instr_rt_idx__T_22_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_22_addr] <= queue_bits_wb_instr_rt_idx__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_23_en & queue_bits_wb_instr_rt_idx__T_23_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_23_addr] <= queue_bits_wb_instr_rt_idx__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_24_en & queue_bits_wb_instr_rt_idx__T_24_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_24_addr] <= queue_bits_wb_instr_rt_idx__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_25_en & queue_bits_wb_instr_rt_idx__T_25_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_25_addr] <= queue_bits_wb_instr_rt_idx__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_26_en & queue_bits_wb_instr_rt_idx__T_26_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_26_addr] <= queue_bits_wb_instr_rt_idx__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_27_en & queue_bits_wb_instr_rt_idx__T_27_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_27_addr] <= queue_bits_wb_instr_rt_idx__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_28_en & queue_bits_wb_instr_rt_idx__T_28_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_28_addr] <= queue_bits_wb_instr_rt_idx__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_29_en & queue_bits_wb_instr_rt_idx__T_29_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_29_addr] <= queue_bits_wb_instr_rt_idx__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_30_en & queue_bits_wb_instr_rt_idx__T_30_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_30_addr] <= queue_bits_wb_instr_rt_idx__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_31_en & queue_bits_wb_instr_rt_idx__T_31_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_31_addr] <= queue_bits_wb_instr_rt_idx__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_32_en & queue_bits_wb_instr_rt_idx__T_32_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_32_addr] <= queue_bits_wb_instr_rt_idx__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_33_en & queue_bits_wb_instr_rt_idx__T_33_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_33_addr] <= queue_bits_wb_instr_rt_idx__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_34_en & queue_bits_wb_instr_rt_idx__T_34_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_34_addr] <= queue_bits_wb_instr_rt_idx__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_35_en & queue_bits_wb_instr_rt_idx__T_35_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_35_addr] <= queue_bits_wb_instr_rt_idx__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_36_en & queue_bits_wb_instr_rt_idx__T_36_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_36_addr] <= queue_bits_wb_instr_rt_idx__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_37_en & queue_bits_wb_instr_rt_idx__T_37_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_37_addr] <= queue_bits_wb_instr_rt_idx__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_38_en & queue_bits_wb_instr_rt_idx__T_38_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_38_addr] <= queue_bits_wb_instr_rt_idx__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_39_en & queue_bits_wb_instr_rt_idx__T_39_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_39_addr] <= queue_bits_wb_instr_rt_idx__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_40_en & queue_bits_wb_instr_rt_idx__T_40_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_40_addr] <= queue_bits_wb_instr_rt_idx__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_41_en & queue_bits_wb_instr_rt_idx__T_41_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_41_addr] <= queue_bits_wb_instr_rt_idx__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_42_en & queue_bits_wb_instr_rt_idx__T_42_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_42_addr] <= queue_bits_wb_instr_rt_idx__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_43_en & queue_bits_wb_instr_rt_idx__T_43_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_43_addr] <= queue_bits_wb_instr_rt_idx__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_44_en & queue_bits_wb_instr_rt_idx__T_44_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_44_addr] <= queue_bits_wb_instr_rt_idx__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_45_en & queue_bits_wb_instr_rt_idx__T_45_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_45_addr] <= queue_bits_wb_instr_rt_idx__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_46_en & queue_bits_wb_instr_rt_idx__T_46_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_46_addr] <= queue_bits_wb_instr_rt_idx__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_47_en & queue_bits_wb_instr_rt_idx__T_47_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_47_addr] <= queue_bits_wb_instr_rt_idx__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_48_en & queue_bits_wb_instr_rt_idx__T_48_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_48_addr] <= queue_bits_wb_instr_rt_idx__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_49_en & queue_bits_wb_instr_rt_idx__T_49_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_49_addr] <= queue_bits_wb_instr_rt_idx__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_50_en & queue_bits_wb_instr_rt_idx__T_50_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_50_addr] <= queue_bits_wb_instr_rt_idx__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_51_en & queue_bits_wb_instr_rt_idx__T_51_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_51_addr] <= queue_bits_wb_instr_rt_idx__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_52_en & queue_bits_wb_instr_rt_idx__T_52_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_52_addr] <= queue_bits_wb_instr_rt_idx__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_53_en & queue_bits_wb_instr_rt_idx__T_53_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_53_addr] <= queue_bits_wb_instr_rt_idx__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_54_en & queue_bits_wb_instr_rt_idx__T_54_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_54_addr] <= queue_bits_wb_instr_rt_idx__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_55_en & queue_bits_wb_instr_rt_idx__T_55_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_55_addr] <= queue_bits_wb_instr_rt_idx__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_56_en & queue_bits_wb_instr_rt_idx__T_56_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_56_addr] <= queue_bits_wb_instr_rt_idx__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_57_en & queue_bits_wb_instr_rt_idx__T_57_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_57_addr] <= queue_bits_wb_instr_rt_idx__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_58_en & queue_bits_wb_instr_rt_idx__T_58_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_58_addr] <= queue_bits_wb_instr_rt_idx__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_59_en & queue_bits_wb_instr_rt_idx__T_59_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_59_addr] <= queue_bits_wb_instr_rt_idx__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_60_en & queue_bits_wb_instr_rt_idx__T_60_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_60_addr] <= queue_bits_wb_instr_rt_idx__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_61_en & queue_bits_wb_instr_rt_idx__T_61_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_61_addr] <= queue_bits_wb_instr_rt_idx__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_62_en & queue_bits_wb_instr_rt_idx__T_62_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_62_addr] <= queue_bits_wb_instr_rt_idx__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_63_en & queue_bits_wb_instr_rt_idx__T_63_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_63_addr] <= queue_bits_wb_instr_rt_idx__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_64_en & queue_bits_wb_instr_rt_idx__T_64_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_64_addr] <= queue_bits_wb_instr_rt_idx__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_65_en & queue_bits_wb_instr_rt_idx__T_65_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_65_addr] <= queue_bits_wb_instr_rt_idx__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_66_en & queue_bits_wb_instr_rt_idx__T_66_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_66_addr] <= queue_bits_wb_instr_rt_idx__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_67_en & queue_bits_wb_instr_rt_idx__T_67_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_67_addr] <= queue_bits_wb_instr_rt_idx__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_68_en & queue_bits_wb_instr_rt_idx__T_68_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_68_addr] <= queue_bits_wb_instr_rt_idx__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_70_en & queue_bits_wb_instr_rt_idx__T_70_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_70_addr] <= queue_bits_wb_instr_rt_idx__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_71_en & queue_bits_wb_instr_rt_idx__T_71_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_71_addr] <= queue_bits_wb_instr_rt_idx__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_72_en & queue_bits_wb_instr_rt_idx__T_72_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_72_addr] <= queue_bits_wb_instr_rt_idx__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_73_en & queue_bits_wb_instr_rt_idx__T_73_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_73_addr] <= queue_bits_wb_instr_rt_idx__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_74_en & queue_bits_wb_instr_rt_idx__T_74_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_74_addr] <= queue_bits_wb_instr_rt_idx__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_75_en & queue_bits_wb_instr_rt_idx__T_75_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_75_addr] <= queue_bits_wb_instr_rt_idx__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_76_en & queue_bits_wb_instr_rt_idx__T_76_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_76_addr] <= queue_bits_wb_instr_rt_idx__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_77_en & queue_bits_wb_instr_rt_idx__T_77_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_77_addr] <= queue_bits_wb_instr_rt_idx__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_78_en & queue_bits_wb_instr_rt_idx__T_78_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_78_addr] <= queue_bits_wb_instr_rt_idx__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_79_en & queue_bits_wb_instr_rt_idx__T_79_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_79_addr] <= queue_bits_wb_instr_rt_idx__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_80_en & queue_bits_wb_instr_rt_idx__T_80_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_80_addr] <= queue_bits_wb_instr_rt_idx__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_81_en & queue_bits_wb_instr_rt_idx__T_81_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_81_addr] <= queue_bits_wb_instr_rt_idx__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_82_en & queue_bits_wb_instr_rt_idx__T_82_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_82_addr] <= queue_bits_wb_instr_rt_idx__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_83_en & queue_bits_wb_instr_rt_idx__T_83_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_83_addr] <= queue_bits_wb_instr_rt_idx__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_84_en & queue_bits_wb_instr_rt_idx__T_84_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_84_addr] <= queue_bits_wb_instr_rt_idx__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_85_en & queue_bits_wb_instr_rt_idx__T_85_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_85_addr] <= queue_bits_wb_instr_rt_idx__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_86_en & queue_bits_wb_instr_rt_idx__T_86_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_86_addr] <= queue_bits_wb_instr_rt_idx__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_87_en & queue_bits_wb_instr_rt_idx__T_87_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_87_addr] <= queue_bits_wb_instr_rt_idx__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_88_en & queue_bits_wb_instr_rt_idx__T_88_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_88_addr] <= queue_bits_wb_instr_rt_idx__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_89_en & queue_bits_wb_instr_rt_idx__T_89_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_89_addr] <= queue_bits_wb_instr_rt_idx__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_90_en & queue_bits_wb_instr_rt_idx__T_90_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_90_addr] <= queue_bits_wb_instr_rt_idx__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_91_en & queue_bits_wb_instr_rt_idx__T_91_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_91_addr] <= queue_bits_wb_instr_rt_idx__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_92_en & queue_bits_wb_instr_rt_idx__T_92_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_92_addr] <= queue_bits_wb_instr_rt_idx__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_93_en & queue_bits_wb_instr_rt_idx__T_93_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_93_addr] <= queue_bits_wb_instr_rt_idx__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_94_en & queue_bits_wb_instr_rt_idx__T_94_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_94_addr] <= queue_bits_wb_instr_rt_idx__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_95_en & queue_bits_wb_instr_rt_idx__T_95_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_95_addr] <= queue_bits_wb_instr_rt_idx__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_96_en & queue_bits_wb_instr_rt_idx__T_96_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_96_addr] <= queue_bits_wb_instr_rt_idx__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_97_en & queue_bits_wb_instr_rt_idx__T_97_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_97_addr] <= queue_bits_wb_instr_rt_idx__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_98_en & queue_bits_wb_instr_rt_idx__T_98_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_98_addr] <= queue_bits_wb_instr_rt_idx__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_99_en & queue_bits_wb_instr_rt_idx__T_99_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_99_addr] <= queue_bits_wb_instr_rt_idx__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_100_en & queue_bits_wb_instr_rt_idx__T_100_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_100_addr] <= queue_bits_wb_instr_rt_idx__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_101_en & queue_bits_wb_instr_rt_idx__T_101_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_101_addr] <= queue_bits_wb_instr_rt_idx__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_102_en & queue_bits_wb_instr_rt_idx__T_102_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_102_addr] <= queue_bits_wb_instr_rt_idx__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_103_en & queue_bits_wb_instr_rt_idx__T_103_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_103_addr] <= queue_bits_wb_instr_rt_idx__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_104_en & queue_bits_wb_instr_rt_idx__T_104_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_104_addr] <= queue_bits_wb_instr_rt_idx__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_105_en & queue_bits_wb_instr_rt_idx__T_105_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_105_addr] <= queue_bits_wb_instr_rt_idx__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_106_en & queue_bits_wb_instr_rt_idx__T_106_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_106_addr] <= queue_bits_wb_instr_rt_idx__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_107_en & queue_bits_wb_instr_rt_idx__T_107_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_107_addr] <= queue_bits_wb_instr_rt_idx__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_108_en & queue_bits_wb_instr_rt_idx__T_108_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_108_addr] <= queue_bits_wb_instr_rt_idx__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_109_en & queue_bits_wb_instr_rt_idx__T_109_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_109_addr] <= queue_bits_wb_instr_rt_idx__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_110_en & queue_bits_wb_instr_rt_idx__T_110_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_110_addr] <= queue_bits_wb_instr_rt_idx__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_111_en & queue_bits_wb_instr_rt_idx__T_111_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_111_addr] <= queue_bits_wb_instr_rt_idx__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_112_en & queue_bits_wb_instr_rt_idx__T_112_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_112_addr] <= queue_bits_wb_instr_rt_idx__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_113_en & queue_bits_wb_instr_rt_idx__T_113_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_113_addr] <= queue_bits_wb_instr_rt_idx__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_114_en & queue_bits_wb_instr_rt_idx__T_114_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_114_addr] <= queue_bits_wb_instr_rt_idx__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_115_en & queue_bits_wb_instr_rt_idx__T_115_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_115_addr] <= queue_bits_wb_instr_rt_idx__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_116_en & queue_bits_wb_instr_rt_idx__T_116_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_116_addr] <= queue_bits_wb_instr_rt_idx__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_117_en & queue_bits_wb_instr_rt_idx__T_117_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_117_addr] <= queue_bits_wb_instr_rt_idx__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_118_en & queue_bits_wb_instr_rt_idx__T_118_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_118_addr] <= queue_bits_wb_instr_rt_idx__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_119_en & queue_bits_wb_instr_rt_idx__T_119_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_119_addr] <= queue_bits_wb_instr_rt_idx__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_120_en & queue_bits_wb_instr_rt_idx__T_120_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_120_addr] <= queue_bits_wb_instr_rt_idx__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_121_en & queue_bits_wb_instr_rt_idx__T_121_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_121_addr] <= queue_bits_wb_instr_rt_idx__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_122_en & queue_bits_wb_instr_rt_idx__T_122_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_122_addr] <= queue_bits_wb_instr_rt_idx__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_123_en & queue_bits_wb_instr_rt_idx__T_123_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_123_addr] <= queue_bits_wb_instr_rt_idx__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_124_en & queue_bits_wb_instr_rt_idx__T_124_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_124_addr] <= queue_bits_wb_instr_rt_idx__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_125_en & queue_bits_wb_instr_rt_idx__T_125_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_125_addr] <= queue_bits_wb_instr_rt_idx__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_126_en & queue_bits_wb_instr_rt_idx__T_126_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_126_addr] <= queue_bits_wb_instr_rt_idx__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_127_en & queue_bits_wb_instr_rt_idx__T_127_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_127_addr] <= queue_bits_wb_instr_rt_idx__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_128_en & queue_bits_wb_instr_rt_idx__T_128_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_128_addr] <= queue_bits_wb_instr_rt_idx__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_129_en & queue_bits_wb_instr_rt_idx__T_129_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_129_addr] <= queue_bits_wb_instr_rt_idx__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_130_en & queue_bits_wb_instr_rt_idx__T_130_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_130_addr] <= queue_bits_wb_instr_rt_idx__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_131_en & queue_bits_wb_instr_rt_idx__T_131_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_131_addr] <= queue_bits_wb_instr_rt_idx__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_132_en & queue_bits_wb_instr_rt_idx__T_132_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_132_addr] <= queue_bits_wb_instr_rt_idx__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx__T_133_en & queue_bits_wb_instr_rt_idx__T_133_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx__T_133_addr] <= queue_bits_wb_instr_rt_idx__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rt_idx_q_head_w_en & queue_bits_wb_instr_rt_idx_q_head_w_mask) begin
      queue_bits_wb_instr_rt_idx[queue_bits_wb_instr_rt_idx_q_head_w_addr] <= queue_bits_wb_instr_rt_idx_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_3_en & queue_bits_wb_instr_rd_idx__T_3_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_3_addr] <= queue_bits_wb_instr_rd_idx__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_4_en & queue_bits_wb_instr_rd_idx__T_4_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_4_addr] <= queue_bits_wb_instr_rd_idx__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_5_en & queue_bits_wb_instr_rd_idx__T_5_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_5_addr] <= queue_bits_wb_instr_rd_idx__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_6_en & queue_bits_wb_instr_rd_idx__T_6_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_6_addr] <= queue_bits_wb_instr_rd_idx__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_7_en & queue_bits_wb_instr_rd_idx__T_7_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_7_addr] <= queue_bits_wb_instr_rd_idx__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_8_en & queue_bits_wb_instr_rd_idx__T_8_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_8_addr] <= queue_bits_wb_instr_rd_idx__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_9_en & queue_bits_wb_instr_rd_idx__T_9_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_9_addr] <= queue_bits_wb_instr_rd_idx__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_10_en & queue_bits_wb_instr_rd_idx__T_10_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_10_addr] <= queue_bits_wb_instr_rd_idx__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_11_en & queue_bits_wb_instr_rd_idx__T_11_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_11_addr] <= queue_bits_wb_instr_rd_idx__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_12_en & queue_bits_wb_instr_rd_idx__T_12_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_12_addr] <= queue_bits_wb_instr_rd_idx__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_13_en & queue_bits_wb_instr_rd_idx__T_13_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_13_addr] <= queue_bits_wb_instr_rd_idx__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_14_en & queue_bits_wb_instr_rd_idx__T_14_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_14_addr] <= queue_bits_wb_instr_rd_idx__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_15_en & queue_bits_wb_instr_rd_idx__T_15_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_15_addr] <= queue_bits_wb_instr_rd_idx__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_16_en & queue_bits_wb_instr_rd_idx__T_16_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_16_addr] <= queue_bits_wb_instr_rd_idx__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_17_en & queue_bits_wb_instr_rd_idx__T_17_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_17_addr] <= queue_bits_wb_instr_rd_idx__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_18_en & queue_bits_wb_instr_rd_idx__T_18_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_18_addr] <= queue_bits_wb_instr_rd_idx__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_19_en & queue_bits_wb_instr_rd_idx__T_19_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_19_addr] <= queue_bits_wb_instr_rd_idx__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_20_en & queue_bits_wb_instr_rd_idx__T_20_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_20_addr] <= queue_bits_wb_instr_rd_idx__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_21_en & queue_bits_wb_instr_rd_idx__T_21_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_21_addr] <= queue_bits_wb_instr_rd_idx__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_22_en & queue_bits_wb_instr_rd_idx__T_22_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_22_addr] <= queue_bits_wb_instr_rd_idx__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_23_en & queue_bits_wb_instr_rd_idx__T_23_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_23_addr] <= queue_bits_wb_instr_rd_idx__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_24_en & queue_bits_wb_instr_rd_idx__T_24_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_24_addr] <= queue_bits_wb_instr_rd_idx__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_25_en & queue_bits_wb_instr_rd_idx__T_25_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_25_addr] <= queue_bits_wb_instr_rd_idx__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_26_en & queue_bits_wb_instr_rd_idx__T_26_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_26_addr] <= queue_bits_wb_instr_rd_idx__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_27_en & queue_bits_wb_instr_rd_idx__T_27_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_27_addr] <= queue_bits_wb_instr_rd_idx__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_28_en & queue_bits_wb_instr_rd_idx__T_28_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_28_addr] <= queue_bits_wb_instr_rd_idx__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_29_en & queue_bits_wb_instr_rd_idx__T_29_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_29_addr] <= queue_bits_wb_instr_rd_idx__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_30_en & queue_bits_wb_instr_rd_idx__T_30_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_30_addr] <= queue_bits_wb_instr_rd_idx__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_31_en & queue_bits_wb_instr_rd_idx__T_31_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_31_addr] <= queue_bits_wb_instr_rd_idx__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_32_en & queue_bits_wb_instr_rd_idx__T_32_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_32_addr] <= queue_bits_wb_instr_rd_idx__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_33_en & queue_bits_wb_instr_rd_idx__T_33_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_33_addr] <= queue_bits_wb_instr_rd_idx__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_34_en & queue_bits_wb_instr_rd_idx__T_34_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_34_addr] <= queue_bits_wb_instr_rd_idx__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_35_en & queue_bits_wb_instr_rd_idx__T_35_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_35_addr] <= queue_bits_wb_instr_rd_idx__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_36_en & queue_bits_wb_instr_rd_idx__T_36_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_36_addr] <= queue_bits_wb_instr_rd_idx__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_37_en & queue_bits_wb_instr_rd_idx__T_37_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_37_addr] <= queue_bits_wb_instr_rd_idx__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_38_en & queue_bits_wb_instr_rd_idx__T_38_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_38_addr] <= queue_bits_wb_instr_rd_idx__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_39_en & queue_bits_wb_instr_rd_idx__T_39_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_39_addr] <= queue_bits_wb_instr_rd_idx__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_40_en & queue_bits_wb_instr_rd_idx__T_40_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_40_addr] <= queue_bits_wb_instr_rd_idx__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_41_en & queue_bits_wb_instr_rd_idx__T_41_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_41_addr] <= queue_bits_wb_instr_rd_idx__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_42_en & queue_bits_wb_instr_rd_idx__T_42_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_42_addr] <= queue_bits_wb_instr_rd_idx__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_43_en & queue_bits_wb_instr_rd_idx__T_43_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_43_addr] <= queue_bits_wb_instr_rd_idx__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_44_en & queue_bits_wb_instr_rd_idx__T_44_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_44_addr] <= queue_bits_wb_instr_rd_idx__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_45_en & queue_bits_wb_instr_rd_idx__T_45_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_45_addr] <= queue_bits_wb_instr_rd_idx__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_46_en & queue_bits_wb_instr_rd_idx__T_46_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_46_addr] <= queue_bits_wb_instr_rd_idx__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_47_en & queue_bits_wb_instr_rd_idx__T_47_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_47_addr] <= queue_bits_wb_instr_rd_idx__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_48_en & queue_bits_wb_instr_rd_idx__T_48_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_48_addr] <= queue_bits_wb_instr_rd_idx__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_49_en & queue_bits_wb_instr_rd_idx__T_49_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_49_addr] <= queue_bits_wb_instr_rd_idx__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_50_en & queue_bits_wb_instr_rd_idx__T_50_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_50_addr] <= queue_bits_wb_instr_rd_idx__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_51_en & queue_bits_wb_instr_rd_idx__T_51_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_51_addr] <= queue_bits_wb_instr_rd_idx__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_52_en & queue_bits_wb_instr_rd_idx__T_52_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_52_addr] <= queue_bits_wb_instr_rd_idx__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_53_en & queue_bits_wb_instr_rd_idx__T_53_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_53_addr] <= queue_bits_wb_instr_rd_idx__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_54_en & queue_bits_wb_instr_rd_idx__T_54_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_54_addr] <= queue_bits_wb_instr_rd_idx__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_55_en & queue_bits_wb_instr_rd_idx__T_55_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_55_addr] <= queue_bits_wb_instr_rd_idx__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_56_en & queue_bits_wb_instr_rd_idx__T_56_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_56_addr] <= queue_bits_wb_instr_rd_idx__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_57_en & queue_bits_wb_instr_rd_idx__T_57_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_57_addr] <= queue_bits_wb_instr_rd_idx__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_58_en & queue_bits_wb_instr_rd_idx__T_58_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_58_addr] <= queue_bits_wb_instr_rd_idx__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_59_en & queue_bits_wb_instr_rd_idx__T_59_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_59_addr] <= queue_bits_wb_instr_rd_idx__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_60_en & queue_bits_wb_instr_rd_idx__T_60_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_60_addr] <= queue_bits_wb_instr_rd_idx__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_61_en & queue_bits_wb_instr_rd_idx__T_61_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_61_addr] <= queue_bits_wb_instr_rd_idx__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_62_en & queue_bits_wb_instr_rd_idx__T_62_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_62_addr] <= queue_bits_wb_instr_rd_idx__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_63_en & queue_bits_wb_instr_rd_idx__T_63_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_63_addr] <= queue_bits_wb_instr_rd_idx__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_64_en & queue_bits_wb_instr_rd_idx__T_64_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_64_addr] <= queue_bits_wb_instr_rd_idx__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_65_en & queue_bits_wb_instr_rd_idx__T_65_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_65_addr] <= queue_bits_wb_instr_rd_idx__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_66_en & queue_bits_wb_instr_rd_idx__T_66_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_66_addr] <= queue_bits_wb_instr_rd_idx__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_67_en & queue_bits_wb_instr_rd_idx__T_67_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_67_addr] <= queue_bits_wb_instr_rd_idx__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_68_en & queue_bits_wb_instr_rd_idx__T_68_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_68_addr] <= queue_bits_wb_instr_rd_idx__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_70_en & queue_bits_wb_instr_rd_idx__T_70_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_70_addr] <= queue_bits_wb_instr_rd_idx__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_71_en & queue_bits_wb_instr_rd_idx__T_71_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_71_addr] <= queue_bits_wb_instr_rd_idx__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_72_en & queue_bits_wb_instr_rd_idx__T_72_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_72_addr] <= queue_bits_wb_instr_rd_idx__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_73_en & queue_bits_wb_instr_rd_idx__T_73_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_73_addr] <= queue_bits_wb_instr_rd_idx__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_74_en & queue_bits_wb_instr_rd_idx__T_74_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_74_addr] <= queue_bits_wb_instr_rd_idx__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_75_en & queue_bits_wb_instr_rd_idx__T_75_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_75_addr] <= queue_bits_wb_instr_rd_idx__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_76_en & queue_bits_wb_instr_rd_idx__T_76_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_76_addr] <= queue_bits_wb_instr_rd_idx__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_77_en & queue_bits_wb_instr_rd_idx__T_77_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_77_addr] <= queue_bits_wb_instr_rd_idx__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_78_en & queue_bits_wb_instr_rd_idx__T_78_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_78_addr] <= queue_bits_wb_instr_rd_idx__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_79_en & queue_bits_wb_instr_rd_idx__T_79_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_79_addr] <= queue_bits_wb_instr_rd_idx__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_80_en & queue_bits_wb_instr_rd_idx__T_80_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_80_addr] <= queue_bits_wb_instr_rd_idx__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_81_en & queue_bits_wb_instr_rd_idx__T_81_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_81_addr] <= queue_bits_wb_instr_rd_idx__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_82_en & queue_bits_wb_instr_rd_idx__T_82_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_82_addr] <= queue_bits_wb_instr_rd_idx__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_83_en & queue_bits_wb_instr_rd_idx__T_83_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_83_addr] <= queue_bits_wb_instr_rd_idx__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_84_en & queue_bits_wb_instr_rd_idx__T_84_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_84_addr] <= queue_bits_wb_instr_rd_idx__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_85_en & queue_bits_wb_instr_rd_idx__T_85_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_85_addr] <= queue_bits_wb_instr_rd_idx__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_86_en & queue_bits_wb_instr_rd_idx__T_86_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_86_addr] <= queue_bits_wb_instr_rd_idx__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_87_en & queue_bits_wb_instr_rd_idx__T_87_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_87_addr] <= queue_bits_wb_instr_rd_idx__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_88_en & queue_bits_wb_instr_rd_idx__T_88_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_88_addr] <= queue_bits_wb_instr_rd_idx__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_89_en & queue_bits_wb_instr_rd_idx__T_89_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_89_addr] <= queue_bits_wb_instr_rd_idx__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_90_en & queue_bits_wb_instr_rd_idx__T_90_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_90_addr] <= queue_bits_wb_instr_rd_idx__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_91_en & queue_bits_wb_instr_rd_idx__T_91_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_91_addr] <= queue_bits_wb_instr_rd_idx__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_92_en & queue_bits_wb_instr_rd_idx__T_92_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_92_addr] <= queue_bits_wb_instr_rd_idx__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_93_en & queue_bits_wb_instr_rd_idx__T_93_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_93_addr] <= queue_bits_wb_instr_rd_idx__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_94_en & queue_bits_wb_instr_rd_idx__T_94_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_94_addr] <= queue_bits_wb_instr_rd_idx__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_95_en & queue_bits_wb_instr_rd_idx__T_95_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_95_addr] <= queue_bits_wb_instr_rd_idx__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_96_en & queue_bits_wb_instr_rd_idx__T_96_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_96_addr] <= queue_bits_wb_instr_rd_idx__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_97_en & queue_bits_wb_instr_rd_idx__T_97_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_97_addr] <= queue_bits_wb_instr_rd_idx__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_98_en & queue_bits_wb_instr_rd_idx__T_98_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_98_addr] <= queue_bits_wb_instr_rd_idx__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_99_en & queue_bits_wb_instr_rd_idx__T_99_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_99_addr] <= queue_bits_wb_instr_rd_idx__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_100_en & queue_bits_wb_instr_rd_idx__T_100_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_100_addr] <= queue_bits_wb_instr_rd_idx__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_101_en & queue_bits_wb_instr_rd_idx__T_101_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_101_addr] <= queue_bits_wb_instr_rd_idx__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_102_en & queue_bits_wb_instr_rd_idx__T_102_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_102_addr] <= queue_bits_wb_instr_rd_idx__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_103_en & queue_bits_wb_instr_rd_idx__T_103_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_103_addr] <= queue_bits_wb_instr_rd_idx__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_104_en & queue_bits_wb_instr_rd_idx__T_104_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_104_addr] <= queue_bits_wb_instr_rd_idx__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_105_en & queue_bits_wb_instr_rd_idx__T_105_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_105_addr] <= queue_bits_wb_instr_rd_idx__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_106_en & queue_bits_wb_instr_rd_idx__T_106_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_106_addr] <= queue_bits_wb_instr_rd_idx__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_107_en & queue_bits_wb_instr_rd_idx__T_107_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_107_addr] <= queue_bits_wb_instr_rd_idx__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_108_en & queue_bits_wb_instr_rd_idx__T_108_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_108_addr] <= queue_bits_wb_instr_rd_idx__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_109_en & queue_bits_wb_instr_rd_idx__T_109_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_109_addr] <= queue_bits_wb_instr_rd_idx__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_110_en & queue_bits_wb_instr_rd_idx__T_110_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_110_addr] <= queue_bits_wb_instr_rd_idx__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_111_en & queue_bits_wb_instr_rd_idx__T_111_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_111_addr] <= queue_bits_wb_instr_rd_idx__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_112_en & queue_bits_wb_instr_rd_idx__T_112_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_112_addr] <= queue_bits_wb_instr_rd_idx__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_113_en & queue_bits_wb_instr_rd_idx__T_113_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_113_addr] <= queue_bits_wb_instr_rd_idx__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_114_en & queue_bits_wb_instr_rd_idx__T_114_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_114_addr] <= queue_bits_wb_instr_rd_idx__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_115_en & queue_bits_wb_instr_rd_idx__T_115_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_115_addr] <= queue_bits_wb_instr_rd_idx__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_116_en & queue_bits_wb_instr_rd_idx__T_116_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_116_addr] <= queue_bits_wb_instr_rd_idx__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_117_en & queue_bits_wb_instr_rd_idx__T_117_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_117_addr] <= queue_bits_wb_instr_rd_idx__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_118_en & queue_bits_wb_instr_rd_idx__T_118_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_118_addr] <= queue_bits_wb_instr_rd_idx__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_119_en & queue_bits_wb_instr_rd_idx__T_119_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_119_addr] <= queue_bits_wb_instr_rd_idx__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_120_en & queue_bits_wb_instr_rd_idx__T_120_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_120_addr] <= queue_bits_wb_instr_rd_idx__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_121_en & queue_bits_wb_instr_rd_idx__T_121_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_121_addr] <= queue_bits_wb_instr_rd_idx__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_122_en & queue_bits_wb_instr_rd_idx__T_122_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_122_addr] <= queue_bits_wb_instr_rd_idx__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_123_en & queue_bits_wb_instr_rd_idx__T_123_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_123_addr] <= queue_bits_wb_instr_rd_idx__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_124_en & queue_bits_wb_instr_rd_idx__T_124_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_124_addr] <= queue_bits_wb_instr_rd_idx__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_125_en & queue_bits_wb_instr_rd_idx__T_125_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_125_addr] <= queue_bits_wb_instr_rd_idx__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_126_en & queue_bits_wb_instr_rd_idx__T_126_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_126_addr] <= queue_bits_wb_instr_rd_idx__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_127_en & queue_bits_wb_instr_rd_idx__T_127_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_127_addr] <= queue_bits_wb_instr_rd_idx__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_128_en & queue_bits_wb_instr_rd_idx__T_128_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_128_addr] <= queue_bits_wb_instr_rd_idx__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_129_en & queue_bits_wb_instr_rd_idx__T_129_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_129_addr] <= queue_bits_wb_instr_rd_idx__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_130_en & queue_bits_wb_instr_rd_idx__T_130_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_130_addr] <= queue_bits_wb_instr_rd_idx__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_131_en & queue_bits_wb_instr_rd_idx__T_131_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_131_addr] <= queue_bits_wb_instr_rd_idx__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_132_en & queue_bits_wb_instr_rd_idx__T_132_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_132_addr] <= queue_bits_wb_instr_rd_idx__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx__T_133_en & queue_bits_wb_instr_rd_idx__T_133_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx__T_133_addr] <= queue_bits_wb_instr_rd_idx__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_rd_idx_q_head_w_en & queue_bits_wb_instr_rd_idx_q_head_w_mask) begin
      queue_bits_wb_instr_rd_idx[queue_bits_wb_instr_rd_idx_q_head_w_addr] <= queue_bits_wb_instr_rd_idx_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_3_en & queue_bits_wb_instr_shamt__T_3_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_3_addr] <= queue_bits_wb_instr_shamt__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_4_en & queue_bits_wb_instr_shamt__T_4_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_4_addr] <= queue_bits_wb_instr_shamt__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_5_en & queue_bits_wb_instr_shamt__T_5_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_5_addr] <= queue_bits_wb_instr_shamt__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_6_en & queue_bits_wb_instr_shamt__T_6_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_6_addr] <= queue_bits_wb_instr_shamt__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_7_en & queue_bits_wb_instr_shamt__T_7_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_7_addr] <= queue_bits_wb_instr_shamt__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_8_en & queue_bits_wb_instr_shamt__T_8_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_8_addr] <= queue_bits_wb_instr_shamt__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_9_en & queue_bits_wb_instr_shamt__T_9_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_9_addr] <= queue_bits_wb_instr_shamt__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_10_en & queue_bits_wb_instr_shamt__T_10_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_10_addr] <= queue_bits_wb_instr_shamt__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_11_en & queue_bits_wb_instr_shamt__T_11_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_11_addr] <= queue_bits_wb_instr_shamt__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_12_en & queue_bits_wb_instr_shamt__T_12_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_12_addr] <= queue_bits_wb_instr_shamt__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_13_en & queue_bits_wb_instr_shamt__T_13_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_13_addr] <= queue_bits_wb_instr_shamt__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_14_en & queue_bits_wb_instr_shamt__T_14_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_14_addr] <= queue_bits_wb_instr_shamt__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_15_en & queue_bits_wb_instr_shamt__T_15_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_15_addr] <= queue_bits_wb_instr_shamt__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_16_en & queue_bits_wb_instr_shamt__T_16_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_16_addr] <= queue_bits_wb_instr_shamt__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_17_en & queue_bits_wb_instr_shamt__T_17_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_17_addr] <= queue_bits_wb_instr_shamt__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_18_en & queue_bits_wb_instr_shamt__T_18_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_18_addr] <= queue_bits_wb_instr_shamt__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_19_en & queue_bits_wb_instr_shamt__T_19_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_19_addr] <= queue_bits_wb_instr_shamt__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_20_en & queue_bits_wb_instr_shamt__T_20_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_20_addr] <= queue_bits_wb_instr_shamt__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_21_en & queue_bits_wb_instr_shamt__T_21_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_21_addr] <= queue_bits_wb_instr_shamt__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_22_en & queue_bits_wb_instr_shamt__T_22_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_22_addr] <= queue_bits_wb_instr_shamt__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_23_en & queue_bits_wb_instr_shamt__T_23_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_23_addr] <= queue_bits_wb_instr_shamt__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_24_en & queue_bits_wb_instr_shamt__T_24_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_24_addr] <= queue_bits_wb_instr_shamt__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_25_en & queue_bits_wb_instr_shamt__T_25_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_25_addr] <= queue_bits_wb_instr_shamt__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_26_en & queue_bits_wb_instr_shamt__T_26_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_26_addr] <= queue_bits_wb_instr_shamt__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_27_en & queue_bits_wb_instr_shamt__T_27_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_27_addr] <= queue_bits_wb_instr_shamt__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_28_en & queue_bits_wb_instr_shamt__T_28_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_28_addr] <= queue_bits_wb_instr_shamt__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_29_en & queue_bits_wb_instr_shamt__T_29_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_29_addr] <= queue_bits_wb_instr_shamt__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_30_en & queue_bits_wb_instr_shamt__T_30_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_30_addr] <= queue_bits_wb_instr_shamt__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_31_en & queue_bits_wb_instr_shamt__T_31_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_31_addr] <= queue_bits_wb_instr_shamt__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_32_en & queue_bits_wb_instr_shamt__T_32_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_32_addr] <= queue_bits_wb_instr_shamt__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_33_en & queue_bits_wb_instr_shamt__T_33_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_33_addr] <= queue_bits_wb_instr_shamt__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_34_en & queue_bits_wb_instr_shamt__T_34_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_34_addr] <= queue_bits_wb_instr_shamt__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_35_en & queue_bits_wb_instr_shamt__T_35_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_35_addr] <= queue_bits_wb_instr_shamt__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_36_en & queue_bits_wb_instr_shamt__T_36_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_36_addr] <= queue_bits_wb_instr_shamt__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_37_en & queue_bits_wb_instr_shamt__T_37_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_37_addr] <= queue_bits_wb_instr_shamt__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_38_en & queue_bits_wb_instr_shamt__T_38_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_38_addr] <= queue_bits_wb_instr_shamt__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_39_en & queue_bits_wb_instr_shamt__T_39_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_39_addr] <= queue_bits_wb_instr_shamt__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_40_en & queue_bits_wb_instr_shamt__T_40_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_40_addr] <= queue_bits_wb_instr_shamt__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_41_en & queue_bits_wb_instr_shamt__T_41_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_41_addr] <= queue_bits_wb_instr_shamt__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_42_en & queue_bits_wb_instr_shamt__T_42_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_42_addr] <= queue_bits_wb_instr_shamt__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_43_en & queue_bits_wb_instr_shamt__T_43_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_43_addr] <= queue_bits_wb_instr_shamt__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_44_en & queue_bits_wb_instr_shamt__T_44_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_44_addr] <= queue_bits_wb_instr_shamt__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_45_en & queue_bits_wb_instr_shamt__T_45_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_45_addr] <= queue_bits_wb_instr_shamt__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_46_en & queue_bits_wb_instr_shamt__T_46_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_46_addr] <= queue_bits_wb_instr_shamt__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_47_en & queue_bits_wb_instr_shamt__T_47_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_47_addr] <= queue_bits_wb_instr_shamt__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_48_en & queue_bits_wb_instr_shamt__T_48_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_48_addr] <= queue_bits_wb_instr_shamt__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_49_en & queue_bits_wb_instr_shamt__T_49_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_49_addr] <= queue_bits_wb_instr_shamt__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_50_en & queue_bits_wb_instr_shamt__T_50_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_50_addr] <= queue_bits_wb_instr_shamt__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_51_en & queue_bits_wb_instr_shamt__T_51_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_51_addr] <= queue_bits_wb_instr_shamt__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_52_en & queue_bits_wb_instr_shamt__T_52_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_52_addr] <= queue_bits_wb_instr_shamt__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_53_en & queue_bits_wb_instr_shamt__T_53_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_53_addr] <= queue_bits_wb_instr_shamt__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_54_en & queue_bits_wb_instr_shamt__T_54_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_54_addr] <= queue_bits_wb_instr_shamt__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_55_en & queue_bits_wb_instr_shamt__T_55_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_55_addr] <= queue_bits_wb_instr_shamt__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_56_en & queue_bits_wb_instr_shamt__T_56_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_56_addr] <= queue_bits_wb_instr_shamt__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_57_en & queue_bits_wb_instr_shamt__T_57_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_57_addr] <= queue_bits_wb_instr_shamt__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_58_en & queue_bits_wb_instr_shamt__T_58_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_58_addr] <= queue_bits_wb_instr_shamt__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_59_en & queue_bits_wb_instr_shamt__T_59_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_59_addr] <= queue_bits_wb_instr_shamt__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_60_en & queue_bits_wb_instr_shamt__T_60_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_60_addr] <= queue_bits_wb_instr_shamt__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_61_en & queue_bits_wb_instr_shamt__T_61_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_61_addr] <= queue_bits_wb_instr_shamt__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_62_en & queue_bits_wb_instr_shamt__T_62_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_62_addr] <= queue_bits_wb_instr_shamt__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_63_en & queue_bits_wb_instr_shamt__T_63_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_63_addr] <= queue_bits_wb_instr_shamt__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_64_en & queue_bits_wb_instr_shamt__T_64_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_64_addr] <= queue_bits_wb_instr_shamt__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_65_en & queue_bits_wb_instr_shamt__T_65_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_65_addr] <= queue_bits_wb_instr_shamt__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_66_en & queue_bits_wb_instr_shamt__T_66_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_66_addr] <= queue_bits_wb_instr_shamt__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_67_en & queue_bits_wb_instr_shamt__T_67_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_67_addr] <= queue_bits_wb_instr_shamt__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_68_en & queue_bits_wb_instr_shamt__T_68_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_68_addr] <= queue_bits_wb_instr_shamt__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_70_en & queue_bits_wb_instr_shamt__T_70_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_70_addr] <= queue_bits_wb_instr_shamt__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_71_en & queue_bits_wb_instr_shamt__T_71_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_71_addr] <= queue_bits_wb_instr_shamt__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_72_en & queue_bits_wb_instr_shamt__T_72_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_72_addr] <= queue_bits_wb_instr_shamt__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_73_en & queue_bits_wb_instr_shamt__T_73_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_73_addr] <= queue_bits_wb_instr_shamt__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_74_en & queue_bits_wb_instr_shamt__T_74_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_74_addr] <= queue_bits_wb_instr_shamt__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_75_en & queue_bits_wb_instr_shamt__T_75_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_75_addr] <= queue_bits_wb_instr_shamt__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_76_en & queue_bits_wb_instr_shamt__T_76_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_76_addr] <= queue_bits_wb_instr_shamt__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_77_en & queue_bits_wb_instr_shamt__T_77_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_77_addr] <= queue_bits_wb_instr_shamt__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_78_en & queue_bits_wb_instr_shamt__T_78_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_78_addr] <= queue_bits_wb_instr_shamt__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_79_en & queue_bits_wb_instr_shamt__T_79_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_79_addr] <= queue_bits_wb_instr_shamt__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_80_en & queue_bits_wb_instr_shamt__T_80_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_80_addr] <= queue_bits_wb_instr_shamt__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_81_en & queue_bits_wb_instr_shamt__T_81_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_81_addr] <= queue_bits_wb_instr_shamt__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_82_en & queue_bits_wb_instr_shamt__T_82_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_82_addr] <= queue_bits_wb_instr_shamt__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_83_en & queue_bits_wb_instr_shamt__T_83_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_83_addr] <= queue_bits_wb_instr_shamt__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_84_en & queue_bits_wb_instr_shamt__T_84_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_84_addr] <= queue_bits_wb_instr_shamt__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_85_en & queue_bits_wb_instr_shamt__T_85_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_85_addr] <= queue_bits_wb_instr_shamt__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_86_en & queue_bits_wb_instr_shamt__T_86_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_86_addr] <= queue_bits_wb_instr_shamt__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_87_en & queue_bits_wb_instr_shamt__T_87_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_87_addr] <= queue_bits_wb_instr_shamt__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_88_en & queue_bits_wb_instr_shamt__T_88_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_88_addr] <= queue_bits_wb_instr_shamt__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_89_en & queue_bits_wb_instr_shamt__T_89_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_89_addr] <= queue_bits_wb_instr_shamt__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_90_en & queue_bits_wb_instr_shamt__T_90_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_90_addr] <= queue_bits_wb_instr_shamt__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_91_en & queue_bits_wb_instr_shamt__T_91_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_91_addr] <= queue_bits_wb_instr_shamt__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_92_en & queue_bits_wb_instr_shamt__T_92_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_92_addr] <= queue_bits_wb_instr_shamt__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_93_en & queue_bits_wb_instr_shamt__T_93_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_93_addr] <= queue_bits_wb_instr_shamt__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_94_en & queue_bits_wb_instr_shamt__T_94_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_94_addr] <= queue_bits_wb_instr_shamt__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_95_en & queue_bits_wb_instr_shamt__T_95_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_95_addr] <= queue_bits_wb_instr_shamt__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_96_en & queue_bits_wb_instr_shamt__T_96_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_96_addr] <= queue_bits_wb_instr_shamt__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_97_en & queue_bits_wb_instr_shamt__T_97_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_97_addr] <= queue_bits_wb_instr_shamt__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_98_en & queue_bits_wb_instr_shamt__T_98_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_98_addr] <= queue_bits_wb_instr_shamt__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_99_en & queue_bits_wb_instr_shamt__T_99_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_99_addr] <= queue_bits_wb_instr_shamt__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_100_en & queue_bits_wb_instr_shamt__T_100_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_100_addr] <= queue_bits_wb_instr_shamt__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_101_en & queue_bits_wb_instr_shamt__T_101_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_101_addr] <= queue_bits_wb_instr_shamt__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_102_en & queue_bits_wb_instr_shamt__T_102_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_102_addr] <= queue_bits_wb_instr_shamt__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_103_en & queue_bits_wb_instr_shamt__T_103_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_103_addr] <= queue_bits_wb_instr_shamt__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_104_en & queue_bits_wb_instr_shamt__T_104_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_104_addr] <= queue_bits_wb_instr_shamt__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_105_en & queue_bits_wb_instr_shamt__T_105_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_105_addr] <= queue_bits_wb_instr_shamt__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_106_en & queue_bits_wb_instr_shamt__T_106_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_106_addr] <= queue_bits_wb_instr_shamt__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_107_en & queue_bits_wb_instr_shamt__T_107_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_107_addr] <= queue_bits_wb_instr_shamt__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_108_en & queue_bits_wb_instr_shamt__T_108_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_108_addr] <= queue_bits_wb_instr_shamt__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_109_en & queue_bits_wb_instr_shamt__T_109_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_109_addr] <= queue_bits_wb_instr_shamt__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_110_en & queue_bits_wb_instr_shamt__T_110_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_110_addr] <= queue_bits_wb_instr_shamt__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_111_en & queue_bits_wb_instr_shamt__T_111_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_111_addr] <= queue_bits_wb_instr_shamt__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_112_en & queue_bits_wb_instr_shamt__T_112_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_112_addr] <= queue_bits_wb_instr_shamt__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_113_en & queue_bits_wb_instr_shamt__T_113_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_113_addr] <= queue_bits_wb_instr_shamt__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_114_en & queue_bits_wb_instr_shamt__T_114_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_114_addr] <= queue_bits_wb_instr_shamt__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_115_en & queue_bits_wb_instr_shamt__T_115_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_115_addr] <= queue_bits_wb_instr_shamt__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_116_en & queue_bits_wb_instr_shamt__T_116_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_116_addr] <= queue_bits_wb_instr_shamt__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_117_en & queue_bits_wb_instr_shamt__T_117_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_117_addr] <= queue_bits_wb_instr_shamt__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_118_en & queue_bits_wb_instr_shamt__T_118_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_118_addr] <= queue_bits_wb_instr_shamt__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_119_en & queue_bits_wb_instr_shamt__T_119_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_119_addr] <= queue_bits_wb_instr_shamt__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_120_en & queue_bits_wb_instr_shamt__T_120_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_120_addr] <= queue_bits_wb_instr_shamt__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_121_en & queue_bits_wb_instr_shamt__T_121_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_121_addr] <= queue_bits_wb_instr_shamt__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_122_en & queue_bits_wb_instr_shamt__T_122_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_122_addr] <= queue_bits_wb_instr_shamt__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_123_en & queue_bits_wb_instr_shamt__T_123_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_123_addr] <= queue_bits_wb_instr_shamt__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_124_en & queue_bits_wb_instr_shamt__T_124_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_124_addr] <= queue_bits_wb_instr_shamt__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_125_en & queue_bits_wb_instr_shamt__T_125_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_125_addr] <= queue_bits_wb_instr_shamt__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_126_en & queue_bits_wb_instr_shamt__T_126_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_126_addr] <= queue_bits_wb_instr_shamt__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_127_en & queue_bits_wb_instr_shamt__T_127_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_127_addr] <= queue_bits_wb_instr_shamt__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_128_en & queue_bits_wb_instr_shamt__T_128_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_128_addr] <= queue_bits_wb_instr_shamt__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_129_en & queue_bits_wb_instr_shamt__T_129_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_129_addr] <= queue_bits_wb_instr_shamt__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_130_en & queue_bits_wb_instr_shamt__T_130_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_130_addr] <= queue_bits_wb_instr_shamt__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_131_en & queue_bits_wb_instr_shamt__T_131_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_131_addr] <= queue_bits_wb_instr_shamt__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_132_en & queue_bits_wb_instr_shamt__T_132_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_132_addr] <= queue_bits_wb_instr_shamt__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt__T_133_en & queue_bits_wb_instr_shamt__T_133_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt__T_133_addr] <= queue_bits_wb_instr_shamt__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_shamt_q_head_w_en & queue_bits_wb_instr_shamt_q_head_w_mask) begin
      queue_bits_wb_instr_shamt[queue_bits_wb_instr_shamt_q_head_w_addr] <= queue_bits_wb_instr_shamt_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_3_en & queue_bits_wb_instr_func__T_3_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_3_addr] <= queue_bits_wb_instr_func__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_4_en & queue_bits_wb_instr_func__T_4_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_4_addr] <= queue_bits_wb_instr_func__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_5_en & queue_bits_wb_instr_func__T_5_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_5_addr] <= queue_bits_wb_instr_func__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_6_en & queue_bits_wb_instr_func__T_6_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_6_addr] <= queue_bits_wb_instr_func__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_7_en & queue_bits_wb_instr_func__T_7_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_7_addr] <= queue_bits_wb_instr_func__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_8_en & queue_bits_wb_instr_func__T_8_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_8_addr] <= queue_bits_wb_instr_func__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_9_en & queue_bits_wb_instr_func__T_9_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_9_addr] <= queue_bits_wb_instr_func__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_10_en & queue_bits_wb_instr_func__T_10_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_10_addr] <= queue_bits_wb_instr_func__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_11_en & queue_bits_wb_instr_func__T_11_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_11_addr] <= queue_bits_wb_instr_func__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_12_en & queue_bits_wb_instr_func__T_12_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_12_addr] <= queue_bits_wb_instr_func__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_13_en & queue_bits_wb_instr_func__T_13_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_13_addr] <= queue_bits_wb_instr_func__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_14_en & queue_bits_wb_instr_func__T_14_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_14_addr] <= queue_bits_wb_instr_func__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_15_en & queue_bits_wb_instr_func__T_15_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_15_addr] <= queue_bits_wb_instr_func__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_16_en & queue_bits_wb_instr_func__T_16_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_16_addr] <= queue_bits_wb_instr_func__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_17_en & queue_bits_wb_instr_func__T_17_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_17_addr] <= queue_bits_wb_instr_func__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_18_en & queue_bits_wb_instr_func__T_18_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_18_addr] <= queue_bits_wb_instr_func__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_19_en & queue_bits_wb_instr_func__T_19_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_19_addr] <= queue_bits_wb_instr_func__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_20_en & queue_bits_wb_instr_func__T_20_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_20_addr] <= queue_bits_wb_instr_func__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_21_en & queue_bits_wb_instr_func__T_21_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_21_addr] <= queue_bits_wb_instr_func__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_22_en & queue_bits_wb_instr_func__T_22_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_22_addr] <= queue_bits_wb_instr_func__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_23_en & queue_bits_wb_instr_func__T_23_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_23_addr] <= queue_bits_wb_instr_func__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_24_en & queue_bits_wb_instr_func__T_24_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_24_addr] <= queue_bits_wb_instr_func__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_25_en & queue_bits_wb_instr_func__T_25_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_25_addr] <= queue_bits_wb_instr_func__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_26_en & queue_bits_wb_instr_func__T_26_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_26_addr] <= queue_bits_wb_instr_func__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_27_en & queue_bits_wb_instr_func__T_27_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_27_addr] <= queue_bits_wb_instr_func__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_28_en & queue_bits_wb_instr_func__T_28_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_28_addr] <= queue_bits_wb_instr_func__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_29_en & queue_bits_wb_instr_func__T_29_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_29_addr] <= queue_bits_wb_instr_func__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_30_en & queue_bits_wb_instr_func__T_30_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_30_addr] <= queue_bits_wb_instr_func__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_31_en & queue_bits_wb_instr_func__T_31_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_31_addr] <= queue_bits_wb_instr_func__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_32_en & queue_bits_wb_instr_func__T_32_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_32_addr] <= queue_bits_wb_instr_func__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_33_en & queue_bits_wb_instr_func__T_33_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_33_addr] <= queue_bits_wb_instr_func__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_34_en & queue_bits_wb_instr_func__T_34_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_34_addr] <= queue_bits_wb_instr_func__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_35_en & queue_bits_wb_instr_func__T_35_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_35_addr] <= queue_bits_wb_instr_func__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_36_en & queue_bits_wb_instr_func__T_36_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_36_addr] <= queue_bits_wb_instr_func__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_37_en & queue_bits_wb_instr_func__T_37_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_37_addr] <= queue_bits_wb_instr_func__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_38_en & queue_bits_wb_instr_func__T_38_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_38_addr] <= queue_bits_wb_instr_func__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_39_en & queue_bits_wb_instr_func__T_39_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_39_addr] <= queue_bits_wb_instr_func__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_40_en & queue_bits_wb_instr_func__T_40_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_40_addr] <= queue_bits_wb_instr_func__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_41_en & queue_bits_wb_instr_func__T_41_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_41_addr] <= queue_bits_wb_instr_func__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_42_en & queue_bits_wb_instr_func__T_42_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_42_addr] <= queue_bits_wb_instr_func__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_43_en & queue_bits_wb_instr_func__T_43_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_43_addr] <= queue_bits_wb_instr_func__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_44_en & queue_bits_wb_instr_func__T_44_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_44_addr] <= queue_bits_wb_instr_func__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_45_en & queue_bits_wb_instr_func__T_45_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_45_addr] <= queue_bits_wb_instr_func__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_46_en & queue_bits_wb_instr_func__T_46_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_46_addr] <= queue_bits_wb_instr_func__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_47_en & queue_bits_wb_instr_func__T_47_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_47_addr] <= queue_bits_wb_instr_func__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_48_en & queue_bits_wb_instr_func__T_48_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_48_addr] <= queue_bits_wb_instr_func__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_49_en & queue_bits_wb_instr_func__T_49_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_49_addr] <= queue_bits_wb_instr_func__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_50_en & queue_bits_wb_instr_func__T_50_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_50_addr] <= queue_bits_wb_instr_func__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_51_en & queue_bits_wb_instr_func__T_51_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_51_addr] <= queue_bits_wb_instr_func__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_52_en & queue_bits_wb_instr_func__T_52_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_52_addr] <= queue_bits_wb_instr_func__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_53_en & queue_bits_wb_instr_func__T_53_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_53_addr] <= queue_bits_wb_instr_func__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_54_en & queue_bits_wb_instr_func__T_54_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_54_addr] <= queue_bits_wb_instr_func__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_55_en & queue_bits_wb_instr_func__T_55_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_55_addr] <= queue_bits_wb_instr_func__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_56_en & queue_bits_wb_instr_func__T_56_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_56_addr] <= queue_bits_wb_instr_func__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_57_en & queue_bits_wb_instr_func__T_57_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_57_addr] <= queue_bits_wb_instr_func__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_58_en & queue_bits_wb_instr_func__T_58_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_58_addr] <= queue_bits_wb_instr_func__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_59_en & queue_bits_wb_instr_func__T_59_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_59_addr] <= queue_bits_wb_instr_func__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_60_en & queue_bits_wb_instr_func__T_60_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_60_addr] <= queue_bits_wb_instr_func__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_61_en & queue_bits_wb_instr_func__T_61_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_61_addr] <= queue_bits_wb_instr_func__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_62_en & queue_bits_wb_instr_func__T_62_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_62_addr] <= queue_bits_wb_instr_func__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_63_en & queue_bits_wb_instr_func__T_63_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_63_addr] <= queue_bits_wb_instr_func__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_64_en & queue_bits_wb_instr_func__T_64_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_64_addr] <= queue_bits_wb_instr_func__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_65_en & queue_bits_wb_instr_func__T_65_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_65_addr] <= queue_bits_wb_instr_func__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_66_en & queue_bits_wb_instr_func__T_66_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_66_addr] <= queue_bits_wb_instr_func__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_67_en & queue_bits_wb_instr_func__T_67_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_67_addr] <= queue_bits_wb_instr_func__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_68_en & queue_bits_wb_instr_func__T_68_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_68_addr] <= queue_bits_wb_instr_func__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_70_en & queue_bits_wb_instr_func__T_70_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_70_addr] <= queue_bits_wb_instr_func__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_71_en & queue_bits_wb_instr_func__T_71_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_71_addr] <= queue_bits_wb_instr_func__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_72_en & queue_bits_wb_instr_func__T_72_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_72_addr] <= queue_bits_wb_instr_func__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_73_en & queue_bits_wb_instr_func__T_73_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_73_addr] <= queue_bits_wb_instr_func__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_74_en & queue_bits_wb_instr_func__T_74_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_74_addr] <= queue_bits_wb_instr_func__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_75_en & queue_bits_wb_instr_func__T_75_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_75_addr] <= queue_bits_wb_instr_func__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_76_en & queue_bits_wb_instr_func__T_76_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_76_addr] <= queue_bits_wb_instr_func__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_77_en & queue_bits_wb_instr_func__T_77_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_77_addr] <= queue_bits_wb_instr_func__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_78_en & queue_bits_wb_instr_func__T_78_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_78_addr] <= queue_bits_wb_instr_func__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_79_en & queue_bits_wb_instr_func__T_79_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_79_addr] <= queue_bits_wb_instr_func__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_80_en & queue_bits_wb_instr_func__T_80_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_80_addr] <= queue_bits_wb_instr_func__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_81_en & queue_bits_wb_instr_func__T_81_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_81_addr] <= queue_bits_wb_instr_func__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_82_en & queue_bits_wb_instr_func__T_82_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_82_addr] <= queue_bits_wb_instr_func__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_83_en & queue_bits_wb_instr_func__T_83_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_83_addr] <= queue_bits_wb_instr_func__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_84_en & queue_bits_wb_instr_func__T_84_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_84_addr] <= queue_bits_wb_instr_func__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_85_en & queue_bits_wb_instr_func__T_85_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_85_addr] <= queue_bits_wb_instr_func__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_86_en & queue_bits_wb_instr_func__T_86_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_86_addr] <= queue_bits_wb_instr_func__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_87_en & queue_bits_wb_instr_func__T_87_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_87_addr] <= queue_bits_wb_instr_func__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_88_en & queue_bits_wb_instr_func__T_88_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_88_addr] <= queue_bits_wb_instr_func__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_89_en & queue_bits_wb_instr_func__T_89_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_89_addr] <= queue_bits_wb_instr_func__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_90_en & queue_bits_wb_instr_func__T_90_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_90_addr] <= queue_bits_wb_instr_func__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_91_en & queue_bits_wb_instr_func__T_91_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_91_addr] <= queue_bits_wb_instr_func__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_92_en & queue_bits_wb_instr_func__T_92_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_92_addr] <= queue_bits_wb_instr_func__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_93_en & queue_bits_wb_instr_func__T_93_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_93_addr] <= queue_bits_wb_instr_func__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_94_en & queue_bits_wb_instr_func__T_94_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_94_addr] <= queue_bits_wb_instr_func__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_95_en & queue_bits_wb_instr_func__T_95_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_95_addr] <= queue_bits_wb_instr_func__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_96_en & queue_bits_wb_instr_func__T_96_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_96_addr] <= queue_bits_wb_instr_func__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_97_en & queue_bits_wb_instr_func__T_97_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_97_addr] <= queue_bits_wb_instr_func__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_98_en & queue_bits_wb_instr_func__T_98_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_98_addr] <= queue_bits_wb_instr_func__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_99_en & queue_bits_wb_instr_func__T_99_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_99_addr] <= queue_bits_wb_instr_func__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_100_en & queue_bits_wb_instr_func__T_100_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_100_addr] <= queue_bits_wb_instr_func__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_101_en & queue_bits_wb_instr_func__T_101_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_101_addr] <= queue_bits_wb_instr_func__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_102_en & queue_bits_wb_instr_func__T_102_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_102_addr] <= queue_bits_wb_instr_func__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_103_en & queue_bits_wb_instr_func__T_103_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_103_addr] <= queue_bits_wb_instr_func__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_104_en & queue_bits_wb_instr_func__T_104_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_104_addr] <= queue_bits_wb_instr_func__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_105_en & queue_bits_wb_instr_func__T_105_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_105_addr] <= queue_bits_wb_instr_func__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_106_en & queue_bits_wb_instr_func__T_106_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_106_addr] <= queue_bits_wb_instr_func__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_107_en & queue_bits_wb_instr_func__T_107_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_107_addr] <= queue_bits_wb_instr_func__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_108_en & queue_bits_wb_instr_func__T_108_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_108_addr] <= queue_bits_wb_instr_func__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_109_en & queue_bits_wb_instr_func__T_109_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_109_addr] <= queue_bits_wb_instr_func__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_110_en & queue_bits_wb_instr_func__T_110_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_110_addr] <= queue_bits_wb_instr_func__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_111_en & queue_bits_wb_instr_func__T_111_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_111_addr] <= queue_bits_wb_instr_func__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_112_en & queue_bits_wb_instr_func__T_112_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_112_addr] <= queue_bits_wb_instr_func__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_113_en & queue_bits_wb_instr_func__T_113_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_113_addr] <= queue_bits_wb_instr_func__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_114_en & queue_bits_wb_instr_func__T_114_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_114_addr] <= queue_bits_wb_instr_func__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_115_en & queue_bits_wb_instr_func__T_115_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_115_addr] <= queue_bits_wb_instr_func__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_116_en & queue_bits_wb_instr_func__T_116_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_116_addr] <= queue_bits_wb_instr_func__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_117_en & queue_bits_wb_instr_func__T_117_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_117_addr] <= queue_bits_wb_instr_func__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_118_en & queue_bits_wb_instr_func__T_118_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_118_addr] <= queue_bits_wb_instr_func__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_119_en & queue_bits_wb_instr_func__T_119_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_119_addr] <= queue_bits_wb_instr_func__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_120_en & queue_bits_wb_instr_func__T_120_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_120_addr] <= queue_bits_wb_instr_func__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_121_en & queue_bits_wb_instr_func__T_121_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_121_addr] <= queue_bits_wb_instr_func__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_122_en & queue_bits_wb_instr_func__T_122_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_122_addr] <= queue_bits_wb_instr_func__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_123_en & queue_bits_wb_instr_func__T_123_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_123_addr] <= queue_bits_wb_instr_func__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_124_en & queue_bits_wb_instr_func__T_124_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_124_addr] <= queue_bits_wb_instr_func__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_125_en & queue_bits_wb_instr_func__T_125_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_125_addr] <= queue_bits_wb_instr_func__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_126_en & queue_bits_wb_instr_func__T_126_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_126_addr] <= queue_bits_wb_instr_func__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_127_en & queue_bits_wb_instr_func__T_127_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_127_addr] <= queue_bits_wb_instr_func__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_128_en & queue_bits_wb_instr_func__T_128_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_128_addr] <= queue_bits_wb_instr_func__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_129_en & queue_bits_wb_instr_func__T_129_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_129_addr] <= queue_bits_wb_instr_func__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_130_en & queue_bits_wb_instr_func__T_130_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_130_addr] <= queue_bits_wb_instr_func__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_131_en & queue_bits_wb_instr_func__T_131_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_131_addr] <= queue_bits_wb_instr_func__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_132_en & queue_bits_wb_instr_func__T_132_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_132_addr] <= queue_bits_wb_instr_func__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func__T_133_en & queue_bits_wb_instr_func__T_133_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func__T_133_addr] <= queue_bits_wb_instr_func__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_instr_func_q_head_w_en & queue_bits_wb_instr_func_q_head_w_mask) begin
      queue_bits_wb_instr_func[queue_bits_wb_instr_func_q_head_w_addr] <= queue_bits_wb_instr_func_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_3_en & queue_bits_wb_rd_idx__T_3_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_3_addr] <= queue_bits_wb_rd_idx__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_4_en & queue_bits_wb_rd_idx__T_4_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_4_addr] <= queue_bits_wb_rd_idx__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_5_en & queue_bits_wb_rd_idx__T_5_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_5_addr] <= queue_bits_wb_rd_idx__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_6_en & queue_bits_wb_rd_idx__T_6_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_6_addr] <= queue_bits_wb_rd_idx__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_7_en & queue_bits_wb_rd_idx__T_7_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_7_addr] <= queue_bits_wb_rd_idx__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_8_en & queue_bits_wb_rd_idx__T_8_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_8_addr] <= queue_bits_wb_rd_idx__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_9_en & queue_bits_wb_rd_idx__T_9_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_9_addr] <= queue_bits_wb_rd_idx__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_10_en & queue_bits_wb_rd_idx__T_10_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_10_addr] <= queue_bits_wb_rd_idx__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_11_en & queue_bits_wb_rd_idx__T_11_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_11_addr] <= queue_bits_wb_rd_idx__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_12_en & queue_bits_wb_rd_idx__T_12_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_12_addr] <= queue_bits_wb_rd_idx__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_13_en & queue_bits_wb_rd_idx__T_13_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_13_addr] <= queue_bits_wb_rd_idx__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_14_en & queue_bits_wb_rd_idx__T_14_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_14_addr] <= queue_bits_wb_rd_idx__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_15_en & queue_bits_wb_rd_idx__T_15_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_15_addr] <= queue_bits_wb_rd_idx__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_16_en & queue_bits_wb_rd_idx__T_16_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_16_addr] <= queue_bits_wb_rd_idx__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_17_en & queue_bits_wb_rd_idx__T_17_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_17_addr] <= queue_bits_wb_rd_idx__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_18_en & queue_bits_wb_rd_idx__T_18_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_18_addr] <= queue_bits_wb_rd_idx__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_19_en & queue_bits_wb_rd_idx__T_19_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_19_addr] <= queue_bits_wb_rd_idx__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_20_en & queue_bits_wb_rd_idx__T_20_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_20_addr] <= queue_bits_wb_rd_idx__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_21_en & queue_bits_wb_rd_idx__T_21_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_21_addr] <= queue_bits_wb_rd_idx__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_22_en & queue_bits_wb_rd_idx__T_22_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_22_addr] <= queue_bits_wb_rd_idx__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_23_en & queue_bits_wb_rd_idx__T_23_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_23_addr] <= queue_bits_wb_rd_idx__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_24_en & queue_bits_wb_rd_idx__T_24_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_24_addr] <= queue_bits_wb_rd_idx__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_25_en & queue_bits_wb_rd_idx__T_25_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_25_addr] <= queue_bits_wb_rd_idx__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_26_en & queue_bits_wb_rd_idx__T_26_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_26_addr] <= queue_bits_wb_rd_idx__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_27_en & queue_bits_wb_rd_idx__T_27_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_27_addr] <= queue_bits_wb_rd_idx__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_28_en & queue_bits_wb_rd_idx__T_28_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_28_addr] <= queue_bits_wb_rd_idx__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_29_en & queue_bits_wb_rd_idx__T_29_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_29_addr] <= queue_bits_wb_rd_idx__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_30_en & queue_bits_wb_rd_idx__T_30_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_30_addr] <= queue_bits_wb_rd_idx__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_31_en & queue_bits_wb_rd_idx__T_31_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_31_addr] <= queue_bits_wb_rd_idx__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_32_en & queue_bits_wb_rd_idx__T_32_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_32_addr] <= queue_bits_wb_rd_idx__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_33_en & queue_bits_wb_rd_idx__T_33_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_33_addr] <= queue_bits_wb_rd_idx__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_34_en & queue_bits_wb_rd_idx__T_34_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_34_addr] <= queue_bits_wb_rd_idx__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_35_en & queue_bits_wb_rd_idx__T_35_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_35_addr] <= queue_bits_wb_rd_idx__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_36_en & queue_bits_wb_rd_idx__T_36_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_36_addr] <= queue_bits_wb_rd_idx__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_37_en & queue_bits_wb_rd_idx__T_37_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_37_addr] <= queue_bits_wb_rd_idx__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_38_en & queue_bits_wb_rd_idx__T_38_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_38_addr] <= queue_bits_wb_rd_idx__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_39_en & queue_bits_wb_rd_idx__T_39_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_39_addr] <= queue_bits_wb_rd_idx__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_40_en & queue_bits_wb_rd_idx__T_40_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_40_addr] <= queue_bits_wb_rd_idx__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_41_en & queue_bits_wb_rd_idx__T_41_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_41_addr] <= queue_bits_wb_rd_idx__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_42_en & queue_bits_wb_rd_idx__T_42_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_42_addr] <= queue_bits_wb_rd_idx__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_43_en & queue_bits_wb_rd_idx__T_43_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_43_addr] <= queue_bits_wb_rd_idx__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_44_en & queue_bits_wb_rd_idx__T_44_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_44_addr] <= queue_bits_wb_rd_idx__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_45_en & queue_bits_wb_rd_idx__T_45_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_45_addr] <= queue_bits_wb_rd_idx__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_46_en & queue_bits_wb_rd_idx__T_46_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_46_addr] <= queue_bits_wb_rd_idx__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_47_en & queue_bits_wb_rd_idx__T_47_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_47_addr] <= queue_bits_wb_rd_idx__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_48_en & queue_bits_wb_rd_idx__T_48_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_48_addr] <= queue_bits_wb_rd_idx__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_49_en & queue_bits_wb_rd_idx__T_49_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_49_addr] <= queue_bits_wb_rd_idx__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_50_en & queue_bits_wb_rd_idx__T_50_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_50_addr] <= queue_bits_wb_rd_idx__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_51_en & queue_bits_wb_rd_idx__T_51_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_51_addr] <= queue_bits_wb_rd_idx__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_52_en & queue_bits_wb_rd_idx__T_52_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_52_addr] <= queue_bits_wb_rd_idx__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_53_en & queue_bits_wb_rd_idx__T_53_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_53_addr] <= queue_bits_wb_rd_idx__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_54_en & queue_bits_wb_rd_idx__T_54_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_54_addr] <= queue_bits_wb_rd_idx__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_55_en & queue_bits_wb_rd_idx__T_55_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_55_addr] <= queue_bits_wb_rd_idx__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_56_en & queue_bits_wb_rd_idx__T_56_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_56_addr] <= queue_bits_wb_rd_idx__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_57_en & queue_bits_wb_rd_idx__T_57_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_57_addr] <= queue_bits_wb_rd_idx__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_58_en & queue_bits_wb_rd_idx__T_58_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_58_addr] <= queue_bits_wb_rd_idx__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_59_en & queue_bits_wb_rd_idx__T_59_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_59_addr] <= queue_bits_wb_rd_idx__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_60_en & queue_bits_wb_rd_idx__T_60_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_60_addr] <= queue_bits_wb_rd_idx__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_61_en & queue_bits_wb_rd_idx__T_61_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_61_addr] <= queue_bits_wb_rd_idx__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_62_en & queue_bits_wb_rd_idx__T_62_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_62_addr] <= queue_bits_wb_rd_idx__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_63_en & queue_bits_wb_rd_idx__T_63_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_63_addr] <= queue_bits_wb_rd_idx__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_64_en & queue_bits_wb_rd_idx__T_64_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_64_addr] <= queue_bits_wb_rd_idx__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_65_en & queue_bits_wb_rd_idx__T_65_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_65_addr] <= queue_bits_wb_rd_idx__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_66_en & queue_bits_wb_rd_idx__T_66_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_66_addr] <= queue_bits_wb_rd_idx__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_67_en & queue_bits_wb_rd_idx__T_67_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_67_addr] <= queue_bits_wb_rd_idx__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_68_en & queue_bits_wb_rd_idx__T_68_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_68_addr] <= queue_bits_wb_rd_idx__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_70_en & queue_bits_wb_rd_idx__T_70_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_70_addr] <= queue_bits_wb_rd_idx__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_71_en & queue_bits_wb_rd_idx__T_71_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_71_addr] <= queue_bits_wb_rd_idx__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_72_en & queue_bits_wb_rd_idx__T_72_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_72_addr] <= queue_bits_wb_rd_idx__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_73_en & queue_bits_wb_rd_idx__T_73_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_73_addr] <= queue_bits_wb_rd_idx__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_74_en & queue_bits_wb_rd_idx__T_74_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_74_addr] <= queue_bits_wb_rd_idx__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_75_en & queue_bits_wb_rd_idx__T_75_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_75_addr] <= queue_bits_wb_rd_idx__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_76_en & queue_bits_wb_rd_idx__T_76_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_76_addr] <= queue_bits_wb_rd_idx__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_77_en & queue_bits_wb_rd_idx__T_77_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_77_addr] <= queue_bits_wb_rd_idx__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_78_en & queue_bits_wb_rd_idx__T_78_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_78_addr] <= queue_bits_wb_rd_idx__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_79_en & queue_bits_wb_rd_idx__T_79_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_79_addr] <= queue_bits_wb_rd_idx__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_80_en & queue_bits_wb_rd_idx__T_80_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_80_addr] <= queue_bits_wb_rd_idx__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_81_en & queue_bits_wb_rd_idx__T_81_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_81_addr] <= queue_bits_wb_rd_idx__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_82_en & queue_bits_wb_rd_idx__T_82_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_82_addr] <= queue_bits_wb_rd_idx__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_83_en & queue_bits_wb_rd_idx__T_83_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_83_addr] <= queue_bits_wb_rd_idx__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_84_en & queue_bits_wb_rd_idx__T_84_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_84_addr] <= queue_bits_wb_rd_idx__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_85_en & queue_bits_wb_rd_idx__T_85_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_85_addr] <= queue_bits_wb_rd_idx__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_86_en & queue_bits_wb_rd_idx__T_86_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_86_addr] <= queue_bits_wb_rd_idx__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_87_en & queue_bits_wb_rd_idx__T_87_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_87_addr] <= queue_bits_wb_rd_idx__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_88_en & queue_bits_wb_rd_idx__T_88_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_88_addr] <= queue_bits_wb_rd_idx__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_89_en & queue_bits_wb_rd_idx__T_89_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_89_addr] <= queue_bits_wb_rd_idx__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_90_en & queue_bits_wb_rd_idx__T_90_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_90_addr] <= queue_bits_wb_rd_idx__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_91_en & queue_bits_wb_rd_idx__T_91_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_91_addr] <= queue_bits_wb_rd_idx__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_92_en & queue_bits_wb_rd_idx__T_92_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_92_addr] <= queue_bits_wb_rd_idx__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_93_en & queue_bits_wb_rd_idx__T_93_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_93_addr] <= queue_bits_wb_rd_idx__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_94_en & queue_bits_wb_rd_idx__T_94_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_94_addr] <= queue_bits_wb_rd_idx__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_95_en & queue_bits_wb_rd_idx__T_95_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_95_addr] <= queue_bits_wb_rd_idx__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_96_en & queue_bits_wb_rd_idx__T_96_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_96_addr] <= queue_bits_wb_rd_idx__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_97_en & queue_bits_wb_rd_idx__T_97_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_97_addr] <= queue_bits_wb_rd_idx__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_98_en & queue_bits_wb_rd_idx__T_98_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_98_addr] <= queue_bits_wb_rd_idx__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_99_en & queue_bits_wb_rd_idx__T_99_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_99_addr] <= queue_bits_wb_rd_idx__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_100_en & queue_bits_wb_rd_idx__T_100_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_100_addr] <= queue_bits_wb_rd_idx__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_101_en & queue_bits_wb_rd_idx__T_101_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_101_addr] <= queue_bits_wb_rd_idx__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_102_en & queue_bits_wb_rd_idx__T_102_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_102_addr] <= queue_bits_wb_rd_idx__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_103_en & queue_bits_wb_rd_idx__T_103_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_103_addr] <= queue_bits_wb_rd_idx__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_104_en & queue_bits_wb_rd_idx__T_104_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_104_addr] <= queue_bits_wb_rd_idx__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_105_en & queue_bits_wb_rd_idx__T_105_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_105_addr] <= queue_bits_wb_rd_idx__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_106_en & queue_bits_wb_rd_idx__T_106_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_106_addr] <= queue_bits_wb_rd_idx__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_107_en & queue_bits_wb_rd_idx__T_107_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_107_addr] <= queue_bits_wb_rd_idx__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_108_en & queue_bits_wb_rd_idx__T_108_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_108_addr] <= queue_bits_wb_rd_idx__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_109_en & queue_bits_wb_rd_idx__T_109_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_109_addr] <= queue_bits_wb_rd_idx__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_110_en & queue_bits_wb_rd_idx__T_110_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_110_addr] <= queue_bits_wb_rd_idx__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_111_en & queue_bits_wb_rd_idx__T_111_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_111_addr] <= queue_bits_wb_rd_idx__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_112_en & queue_bits_wb_rd_idx__T_112_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_112_addr] <= queue_bits_wb_rd_idx__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_113_en & queue_bits_wb_rd_idx__T_113_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_113_addr] <= queue_bits_wb_rd_idx__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_114_en & queue_bits_wb_rd_idx__T_114_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_114_addr] <= queue_bits_wb_rd_idx__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_115_en & queue_bits_wb_rd_idx__T_115_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_115_addr] <= queue_bits_wb_rd_idx__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_116_en & queue_bits_wb_rd_idx__T_116_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_116_addr] <= queue_bits_wb_rd_idx__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_117_en & queue_bits_wb_rd_idx__T_117_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_117_addr] <= queue_bits_wb_rd_idx__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_118_en & queue_bits_wb_rd_idx__T_118_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_118_addr] <= queue_bits_wb_rd_idx__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_119_en & queue_bits_wb_rd_idx__T_119_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_119_addr] <= queue_bits_wb_rd_idx__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_120_en & queue_bits_wb_rd_idx__T_120_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_120_addr] <= queue_bits_wb_rd_idx__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_121_en & queue_bits_wb_rd_idx__T_121_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_121_addr] <= queue_bits_wb_rd_idx__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_122_en & queue_bits_wb_rd_idx__T_122_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_122_addr] <= queue_bits_wb_rd_idx__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_123_en & queue_bits_wb_rd_idx__T_123_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_123_addr] <= queue_bits_wb_rd_idx__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_124_en & queue_bits_wb_rd_idx__T_124_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_124_addr] <= queue_bits_wb_rd_idx__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_125_en & queue_bits_wb_rd_idx__T_125_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_125_addr] <= queue_bits_wb_rd_idx__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_126_en & queue_bits_wb_rd_idx__T_126_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_126_addr] <= queue_bits_wb_rd_idx__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_127_en & queue_bits_wb_rd_idx__T_127_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_127_addr] <= queue_bits_wb_rd_idx__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_128_en & queue_bits_wb_rd_idx__T_128_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_128_addr] <= queue_bits_wb_rd_idx__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_129_en & queue_bits_wb_rd_idx__T_129_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_129_addr] <= queue_bits_wb_rd_idx__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_130_en & queue_bits_wb_rd_idx__T_130_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_130_addr] <= queue_bits_wb_rd_idx__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_131_en & queue_bits_wb_rd_idx__T_131_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_131_addr] <= queue_bits_wb_rd_idx__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_132_en & queue_bits_wb_rd_idx__T_132_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_132_addr] <= queue_bits_wb_rd_idx__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx__T_133_en & queue_bits_wb_rd_idx__T_133_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx__T_133_addr] <= queue_bits_wb_rd_idx__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_rd_idx_q_head_w_en & queue_bits_wb_rd_idx_q_head_w_mask) begin
      queue_bits_wb_rd_idx[queue_bits_wb_rd_idx_q_head_w_addr] <= queue_bits_wb_rd_idx_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_3_en & queue_bits_wb_ip7__T_3_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_3_addr] <= queue_bits_wb_ip7__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_4_en & queue_bits_wb_ip7__T_4_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_4_addr] <= queue_bits_wb_ip7__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_5_en & queue_bits_wb_ip7__T_5_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_5_addr] <= queue_bits_wb_ip7__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_6_en & queue_bits_wb_ip7__T_6_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_6_addr] <= queue_bits_wb_ip7__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_7_en & queue_bits_wb_ip7__T_7_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_7_addr] <= queue_bits_wb_ip7__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_8_en & queue_bits_wb_ip7__T_8_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_8_addr] <= queue_bits_wb_ip7__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_9_en & queue_bits_wb_ip7__T_9_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_9_addr] <= queue_bits_wb_ip7__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_10_en & queue_bits_wb_ip7__T_10_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_10_addr] <= queue_bits_wb_ip7__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_11_en & queue_bits_wb_ip7__T_11_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_11_addr] <= queue_bits_wb_ip7__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_12_en & queue_bits_wb_ip7__T_12_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_12_addr] <= queue_bits_wb_ip7__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_13_en & queue_bits_wb_ip7__T_13_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_13_addr] <= queue_bits_wb_ip7__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_14_en & queue_bits_wb_ip7__T_14_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_14_addr] <= queue_bits_wb_ip7__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_15_en & queue_bits_wb_ip7__T_15_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_15_addr] <= queue_bits_wb_ip7__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_16_en & queue_bits_wb_ip7__T_16_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_16_addr] <= queue_bits_wb_ip7__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_17_en & queue_bits_wb_ip7__T_17_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_17_addr] <= queue_bits_wb_ip7__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_18_en & queue_bits_wb_ip7__T_18_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_18_addr] <= queue_bits_wb_ip7__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_19_en & queue_bits_wb_ip7__T_19_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_19_addr] <= queue_bits_wb_ip7__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_20_en & queue_bits_wb_ip7__T_20_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_20_addr] <= queue_bits_wb_ip7__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_21_en & queue_bits_wb_ip7__T_21_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_21_addr] <= queue_bits_wb_ip7__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_22_en & queue_bits_wb_ip7__T_22_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_22_addr] <= queue_bits_wb_ip7__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_23_en & queue_bits_wb_ip7__T_23_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_23_addr] <= queue_bits_wb_ip7__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_24_en & queue_bits_wb_ip7__T_24_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_24_addr] <= queue_bits_wb_ip7__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_25_en & queue_bits_wb_ip7__T_25_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_25_addr] <= queue_bits_wb_ip7__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_26_en & queue_bits_wb_ip7__T_26_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_26_addr] <= queue_bits_wb_ip7__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_27_en & queue_bits_wb_ip7__T_27_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_27_addr] <= queue_bits_wb_ip7__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_28_en & queue_bits_wb_ip7__T_28_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_28_addr] <= queue_bits_wb_ip7__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_29_en & queue_bits_wb_ip7__T_29_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_29_addr] <= queue_bits_wb_ip7__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_30_en & queue_bits_wb_ip7__T_30_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_30_addr] <= queue_bits_wb_ip7__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_31_en & queue_bits_wb_ip7__T_31_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_31_addr] <= queue_bits_wb_ip7__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_32_en & queue_bits_wb_ip7__T_32_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_32_addr] <= queue_bits_wb_ip7__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_33_en & queue_bits_wb_ip7__T_33_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_33_addr] <= queue_bits_wb_ip7__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_34_en & queue_bits_wb_ip7__T_34_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_34_addr] <= queue_bits_wb_ip7__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_35_en & queue_bits_wb_ip7__T_35_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_35_addr] <= queue_bits_wb_ip7__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_36_en & queue_bits_wb_ip7__T_36_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_36_addr] <= queue_bits_wb_ip7__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_37_en & queue_bits_wb_ip7__T_37_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_37_addr] <= queue_bits_wb_ip7__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_38_en & queue_bits_wb_ip7__T_38_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_38_addr] <= queue_bits_wb_ip7__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_39_en & queue_bits_wb_ip7__T_39_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_39_addr] <= queue_bits_wb_ip7__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_40_en & queue_bits_wb_ip7__T_40_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_40_addr] <= queue_bits_wb_ip7__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_41_en & queue_bits_wb_ip7__T_41_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_41_addr] <= queue_bits_wb_ip7__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_42_en & queue_bits_wb_ip7__T_42_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_42_addr] <= queue_bits_wb_ip7__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_43_en & queue_bits_wb_ip7__T_43_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_43_addr] <= queue_bits_wb_ip7__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_44_en & queue_bits_wb_ip7__T_44_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_44_addr] <= queue_bits_wb_ip7__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_45_en & queue_bits_wb_ip7__T_45_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_45_addr] <= queue_bits_wb_ip7__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_46_en & queue_bits_wb_ip7__T_46_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_46_addr] <= queue_bits_wb_ip7__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_47_en & queue_bits_wb_ip7__T_47_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_47_addr] <= queue_bits_wb_ip7__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_48_en & queue_bits_wb_ip7__T_48_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_48_addr] <= queue_bits_wb_ip7__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_49_en & queue_bits_wb_ip7__T_49_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_49_addr] <= queue_bits_wb_ip7__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_50_en & queue_bits_wb_ip7__T_50_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_50_addr] <= queue_bits_wb_ip7__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_51_en & queue_bits_wb_ip7__T_51_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_51_addr] <= queue_bits_wb_ip7__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_52_en & queue_bits_wb_ip7__T_52_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_52_addr] <= queue_bits_wb_ip7__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_53_en & queue_bits_wb_ip7__T_53_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_53_addr] <= queue_bits_wb_ip7__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_54_en & queue_bits_wb_ip7__T_54_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_54_addr] <= queue_bits_wb_ip7__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_55_en & queue_bits_wb_ip7__T_55_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_55_addr] <= queue_bits_wb_ip7__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_56_en & queue_bits_wb_ip7__T_56_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_56_addr] <= queue_bits_wb_ip7__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_57_en & queue_bits_wb_ip7__T_57_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_57_addr] <= queue_bits_wb_ip7__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_58_en & queue_bits_wb_ip7__T_58_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_58_addr] <= queue_bits_wb_ip7__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_59_en & queue_bits_wb_ip7__T_59_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_59_addr] <= queue_bits_wb_ip7__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_60_en & queue_bits_wb_ip7__T_60_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_60_addr] <= queue_bits_wb_ip7__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_61_en & queue_bits_wb_ip7__T_61_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_61_addr] <= queue_bits_wb_ip7__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_62_en & queue_bits_wb_ip7__T_62_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_62_addr] <= queue_bits_wb_ip7__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_63_en & queue_bits_wb_ip7__T_63_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_63_addr] <= queue_bits_wb_ip7__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_64_en & queue_bits_wb_ip7__T_64_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_64_addr] <= queue_bits_wb_ip7__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_65_en & queue_bits_wb_ip7__T_65_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_65_addr] <= queue_bits_wb_ip7__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_66_en & queue_bits_wb_ip7__T_66_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_66_addr] <= queue_bits_wb_ip7__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_67_en & queue_bits_wb_ip7__T_67_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_67_addr] <= queue_bits_wb_ip7__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_68_en & queue_bits_wb_ip7__T_68_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_68_addr] <= queue_bits_wb_ip7__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_70_en & queue_bits_wb_ip7__T_70_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_70_addr] <= queue_bits_wb_ip7__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_71_en & queue_bits_wb_ip7__T_71_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_71_addr] <= queue_bits_wb_ip7__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_72_en & queue_bits_wb_ip7__T_72_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_72_addr] <= queue_bits_wb_ip7__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_73_en & queue_bits_wb_ip7__T_73_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_73_addr] <= queue_bits_wb_ip7__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_74_en & queue_bits_wb_ip7__T_74_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_74_addr] <= queue_bits_wb_ip7__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_75_en & queue_bits_wb_ip7__T_75_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_75_addr] <= queue_bits_wb_ip7__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_76_en & queue_bits_wb_ip7__T_76_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_76_addr] <= queue_bits_wb_ip7__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_77_en & queue_bits_wb_ip7__T_77_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_77_addr] <= queue_bits_wb_ip7__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_78_en & queue_bits_wb_ip7__T_78_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_78_addr] <= queue_bits_wb_ip7__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_79_en & queue_bits_wb_ip7__T_79_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_79_addr] <= queue_bits_wb_ip7__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_80_en & queue_bits_wb_ip7__T_80_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_80_addr] <= queue_bits_wb_ip7__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_81_en & queue_bits_wb_ip7__T_81_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_81_addr] <= queue_bits_wb_ip7__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_82_en & queue_bits_wb_ip7__T_82_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_82_addr] <= queue_bits_wb_ip7__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_83_en & queue_bits_wb_ip7__T_83_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_83_addr] <= queue_bits_wb_ip7__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_84_en & queue_bits_wb_ip7__T_84_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_84_addr] <= queue_bits_wb_ip7__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_85_en & queue_bits_wb_ip7__T_85_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_85_addr] <= queue_bits_wb_ip7__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_86_en & queue_bits_wb_ip7__T_86_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_86_addr] <= queue_bits_wb_ip7__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_87_en & queue_bits_wb_ip7__T_87_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_87_addr] <= queue_bits_wb_ip7__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_88_en & queue_bits_wb_ip7__T_88_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_88_addr] <= queue_bits_wb_ip7__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_89_en & queue_bits_wb_ip7__T_89_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_89_addr] <= queue_bits_wb_ip7__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_90_en & queue_bits_wb_ip7__T_90_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_90_addr] <= queue_bits_wb_ip7__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_91_en & queue_bits_wb_ip7__T_91_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_91_addr] <= queue_bits_wb_ip7__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_92_en & queue_bits_wb_ip7__T_92_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_92_addr] <= queue_bits_wb_ip7__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_93_en & queue_bits_wb_ip7__T_93_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_93_addr] <= queue_bits_wb_ip7__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_94_en & queue_bits_wb_ip7__T_94_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_94_addr] <= queue_bits_wb_ip7__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_95_en & queue_bits_wb_ip7__T_95_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_95_addr] <= queue_bits_wb_ip7__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_96_en & queue_bits_wb_ip7__T_96_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_96_addr] <= queue_bits_wb_ip7__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_97_en & queue_bits_wb_ip7__T_97_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_97_addr] <= queue_bits_wb_ip7__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_98_en & queue_bits_wb_ip7__T_98_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_98_addr] <= queue_bits_wb_ip7__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_99_en & queue_bits_wb_ip7__T_99_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_99_addr] <= queue_bits_wb_ip7__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_100_en & queue_bits_wb_ip7__T_100_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_100_addr] <= queue_bits_wb_ip7__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_101_en & queue_bits_wb_ip7__T_101_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_101_addr] <= queue_bits_wb_ip7__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_102_en & queue_bits_wb_ip7__T_102_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_102_addr] <= queue_bits_wb_ip7__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_103_en & queue_bits_wb_ip7__T_103_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_103_addr] <= queue_bits_wb_ip7__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_104_en & queue_bits_wb_ip7__T_104_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_104_addr] <= queue_bits_wb_ip7__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_105_en & queue_bits_wb_ip7__T_105_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_105_addr] <= queue_bits_wb_ip7__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_106_en & queue_bits_wb_ip7__T_106_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_106_addr] <= queue_bits_wb_ip7__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_107_en & queue_bits_wb_ip7__T_107_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_107_addr] <= queue_bits_wb_ip7__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_108_en & queue_bits_wb_ip7__T_108_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_108_addr] <= queue_bits_wb_ip7__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_109_en & queue_bits_wb_ip7__T_109_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_109_addr] <= queue_bits_wb_ip7__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_110_en & queue_bits_wb_ip7__T_110_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_110_addr] <= queue_bits_wb_ip7__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_111_en & queue_bits_wb_ip7__T_111_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_111_addr] <= queue_bits_wb_ip7__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_112_en & queue_bits_wb_ip7__T_112_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_112_addr] <= queue_bits_wb_ip7__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_113_en & queue_bits_wb_ip7__T_113_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_113_addr] <= queue_bits_wb_ip7__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_114_en & queue_bits_wb_ip7__T_114_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_114_addr] <= queue_bits_wb_ip7__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_115_en & queue_bits_wb_ip7__T_115_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_115_addr] <= queue_bits_wb_ip7__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_116_en & queue_bits_wb_ip7__T_116_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_116_addr] <= queue_bits_wb_ip7__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_117_en & queue_bits_wb_ip7__T_117_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_117_addr] <= queue_bits_wb_ip7__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_118_en & queue_bits_wb_ip7__T_118_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_118_addr] <= queue_bits_wb_ip7__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_119_en & queue_bits_wb_ip7__T_119_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_119_addr] <= queue_bits_wb_ip7__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_120_en & queue_bits_wb_ip7__T_120_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_120_addr] <= queue_bits_wb_ip7__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_121_en & queue_bits_wb_ip7__T_121_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_121_addr] <= queue_bits_wb_ip7__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_122_en & queue_bits_wb_ip7__T_122_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_122_addr] <= queue_bits_wb_ip7__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_123_en & queue_bits_wb_ip7__T_123_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_123_addr] <= queue_bits_wb_ip7__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_124_en & queue_bits_wb_ip7__T_124_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_124_addr] <= queue_bits_wb_ip7__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_125_en & queue_bits_wb_ip7__T_125_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_125_addr] <= queue_bits_wb_ip7__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_126_en & queue_bits_wb_ip7__T_126_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_126_addr] <= queue_bits_wb_ip7__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_127_en & queue_bits_wb_ip7__T_127_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_127_addr] <= queue_bits_wb_ip7__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_128_en & queue_bits_wb_ip7__T_128_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_128_addr] <= queue_bits_wb_ip7__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_129_en & queue_bits_wb_ip7__T_129_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_129_addr] <= queue_bits_wb_ip7__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_130_en & queue_bits_wb_ip7__T_130_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_130_addr] <= queue_bits_wb_ip7__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_131_en & queue_bits_wb_ip7__T_131_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_131_addr] <= queue_bits_wb_ip7__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_132_en & queue_bits_wb_ip7__T_132_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_132_addr] <= queue_bits_wb_ip7__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7__T_133_en & queue_bits_wb_ip7__T_133_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7__T_133_addr] <= queue_bits_wb_ip7__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_ip7_q_head_w_en & queue_bits_wb_ip7_q_head_w_mask) begin
      queue_bits_wb_ip7[queue_bits_wb_ip7_q_head_w_addr] <= queue_bits_wb_ip7_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_3_en & queue_bits_wb_is_ds__T_3_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_3_addr] <= queue_bits_wb_is_ds__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_4_en & queue_bits_wb_is_ds__T_4_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_4_addr] <= queue_bits_wb_is_ds__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_5_en & queue_bits_wb_is_ds__T_5_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_5_addr] <= queue_bits_wb_is_ds__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_6_en & queue_bits_wb_is_ds__T_6_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_6_addr] <= queue_bits_wb_is_ds__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_7_en & queue_bits_wb_is_ds__T_7_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_7_addr] <= queue_bits_wb_is_ds__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_8_en & queue_bits_wb_is_ds__T_8_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_8_addr] <= queue_bits_wb_is_ds__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_9_en & queue_bits_wb_is_ds__T_9_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_9_addr] <= queue_bits_wb_is_ds__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_10_en & queue_bits_wb_is_ds__T_10_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_10_addr] <= queue_bits_wb_is_ds__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_11_en & queue_bits_wb_is_ds__T_11_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_11_addr] <= queue_bits_wb_is_ds__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_12_en & queue_bits_wb_is_ds__T_12_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_12_addr] <= queue_bits_wb_is_ds__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_13_en & queue_bits_wb_is_ds__T_13_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_13_addr] <= queue_bits_wb_is_ds__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_14_en & queue_bits_wb_is_ds__T_14_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_14_addr] <= queue_bits_wb_is_ds__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_15_en & queue_bits_wb_is_ds__T_15_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_15_addr] <= queue_bits_wb_is_ds__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_16_en & queue_bits_wb_is_ds__T_16_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_16_addr] <= queue_bits_wb_is_ds__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_17_en & queue_bits_wb_is_ds__T_17_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_17_addr] <= queue_bits_wb_is_ds__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_18_en & queue_bits_wb_is_ds__T_18_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_18_addr] <= queue_bits_wb_is_ds__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_19_en & queue_bits_wb_is_ds__T_19_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_19_addr] <= queue_bits_wb_is_ds__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_20_en & queue_bits_wb_is_ds__T_20_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_20_addr] <= queue_bits_wb_is_ds__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_21_en & queue_bits_wb_is_ds__T_21_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_21_addr] <= queue_bits_wb_is_ds__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_22_en & queue_bits_wb_is_ds__T_22_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_22_addr] <= queue_bits_wb_is_ds__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_23_en & queue_bits_wb_is_ds__T_23_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_23_addr] <= queue_bits_wb_is_ds__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_24_en & queue_bits_wb_is_ds__T_24_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_24_addr] <= queue_bits_wb_is_ds__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_25_en & queue_bits_wb_is_ds__T_25_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_25_addr] <= queue_bits_wb_is_ds__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_26_en & queue_bits_wb_is_ds__T_26_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_26_addr] <= queue_bits_wb_is_ds__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_27_en & queue_bits_wb_is_ds__T_27_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_27_addr] <= queue_bits_wb_is_ds__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_28_en & queue_bits_wb_is_ds__T_28_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_28_addr] <= queue_bits_wb_is_ds__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_29_en & queue_bits_wb_is_ds__T_29_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_29_addr] <= queue_bits_wb_is_ds__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_30_en & queue_bits_wb_is_ds__T_30_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_30_addr] <= queue_bits_wb_is_ds__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_31_en & queue_bits_wb_is_ds__T_31_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_31_addr] <= queue_bits_wb_is_ds__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_32_en & queue_bits_wb_is_ds__T_32_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_32_addr] <= queue_bits_wb_is_ds__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_33_en & queue_bits_wb_is_ds__T_33_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_33_addr] <= queue_bits_wb_is_ds__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_34_en & queue_bits_wb_is_ds__T_34_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_34_addr] <= queue_bits_wb_is_ds__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_35_en & queue_bits_wb_is_ds__T_35_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_35_addr] <= queue_bits_wb_is_ds__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_36_en & queue_bits_wb_is_ds__T_36_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_36_addr] <= queue_bits_wb_is_ds__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_37_en & queue_bits_wb_is_ds__T_37_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_37_addr] <= queue_bits_wb_is_ds__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_38_en & queue_bits_wb_is_ds__T_38_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_38_addr] <= queue_bits_wb_is_ds__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_39_en & queue_bits_wb_is_ds__T_39_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_39_addr] <= queue_bits_wb_is_ds__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_40_en & queue_bits_wb_is_ds__T_40_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_40_addr] <= queue_bits_wb_is_ds__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_41_en & queue_bits_wb_is_ds__T_41_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_41_addr] <= queue_bits_wb_is_ds__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_42_en & queue_bits_wb_is_ds__T_42_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_42_addr] <= queue_bits_wb_is_ds__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_43_en & queue_bits_wb_is_ds__T_43_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_43_addr] <= queue_bits_wb_is_ds__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_44_en & queue_bits_wb_is_ds__T_44_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_44_addr] <= queue_bits_wb_is_ds__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_45_en & queue_bits_wb_is_ds__T_45_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_45_addr] <= queue_bits_wb_is_ds__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_46_en & queue_bits_wb_is_ds__T_46_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_46_addr] <= queue_bits_wb_is_ds__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_47_en & queue_bits_wb_is_ds__T_47_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_47_addr] <= queue_bits_wb_is_ds__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_48_en & queue_bits_wb_is_ds__T_48_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_48_addr] <= queue_bits_wb_is_ds__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_49_en & queue_bits_wb_is_ds__T_49_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_49_addr] <= queue_bits_wb_is_ds__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_50_en & queue_bits_wb_is_ds__T_50_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_50_addr] <= queue_bits_wb_is_ds__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_51_en & queue_bits_wb_is_ds__T_51_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_51_addr] <= queue_bits_wb_is_ds__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_52_en & queue_bits_wb_is_ds__T_52_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_52_addr] <= queue_bits_wb_is_ds__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_53_en & queue_bits_wb_is_ds__T_53_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_53_addr] <= queue_bits_wb_is_ds__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_54_en & queue_bits_wb_is_ds__T_54_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_54_addr] <= queue_bits_wb_is_ds__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_55_en & queue_bits_wb_is_ds__T_55_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_55_addr] <= queue_bits_wb_is_ds__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_56_en & queue_bits_wb_is_ds__T_56_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_56_addr] <= queue_bits_wb_is_ds__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_57_en & queue_bits_wb_is_ds__T_57_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_57_addr] <= queue_bits_wb_is_ds__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_58_en & queue_bits_wb_is_ds__T_58_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_58_addr] <= queue_bits_wb_is_ds__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_59_en & queue_bits_wb_is_ds__T_59_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_59_addr] <= queue_bits_wb_is_ds__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_60_en & queue_bits_wb_is_ds__T_60_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_60_addr] <= queue_bits_wb_is_ds__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_61_en & queue_bits_wb_is_ds__T_61_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_61_addr] <= queue_bits_wb_is_ds__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_62_en & queue_bits_wb_is_ds__T_62_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_62_addr] <= queue_bits_wb_is_ds__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_63_en & queue_bits_wb_is_ds__T_63_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_63_addr] <= queue_bits_wb_is_ds__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_64_en & queue_bits_wb_is_ds__T_64_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_64_addr] <= queue_bits_wb_is_ds__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_65_en & queue_bits_wb_is_ds__T_65_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_65_addr] <= queue_bits_wb_is_ds__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_66_en & queue_bits_wb_is_ds__T_66_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_66_addr] <= queue_bits_wb_is_ds__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_67_en & queue_bits_wb_is_ds__T_67_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_67_addr] <= queue_bits_wb_is_ds__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_68_en & queue_bits_wb_is_ds__T_68_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_68_addr] <= queue_bits_wb_is_ds__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_70_en & queue_bits_wb_is_ds__T_70_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_70_addr] <= queue_bits_wb_is_ds__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_71_en & queue_bits_wb_is_ds__T_71_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_71_addr] <= queue_bits_wb_is_ds__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_72_en & queue_bits_wb_is_ds__T_72_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_72_addr] <= queue_bits_wb_is_ds__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_73_en & queue_bits_wb_is_ds__T_73_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_73_addr] <= queue_bits_wb_is_ds__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_74_en & queue_bits_wb_is_ds__T_74_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_74_addr] <= queue_bits_wb_is_ds__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_75_en & queue_bits_wb_is_ds__T_75_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_75_addr] <= queue_bits_wb_is_ds__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_76_en & queue_bits_wb_is_ds__T_76_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_76_addr] <= queue_bits_wb_is_ds__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_77_en & queue_bits_wb_is_ds__T_77_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_77_addr] <= queue_bits_wb_is_ds__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_78_en & queue_bits_wb_is_ds__T_78_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_78_addr] <= queue_bits_wb_is_ds__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_79_en & queue_bits_wb_is_ds__T_79_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_79_addr] <= queue_bits_wb_is_ds__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_80_en & queue_bits_wb_is_ds__T_80_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_80_addr] <= queue_bits_wb_is_ds__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_81_en & queue_bits_wb_is_ds__T_81_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_81_addr] <= queue_bits_wb_is_ds__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_82_en & queue_bits_wb_is_ds__T_82_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_82_addr] <= queue_bits_wb_is_ds__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_83_en & queue_bits_wb_is_ds__T_83_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_83_addr] <= queue_bits_wb_is_ds__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_84_en & queue_bits_wb_is_ds__T_84_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_84_addr] <= queue_bits_wb_is_ds__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_85_en & queue_bits_wb_is_ds__T_85_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_85_addr] <= queue_bits_wb_is_ds__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_86_en & queue_bits_wb_is_ds__T_86_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_86_addr] <= queue_bits_wb_is_ds__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_87_en & queue_bits_wb_is_ds__T_87_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_87_addr] <= queue_bits_wb_is_ds__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_88_en & queue_bits_wb_is_ds__T_88_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_88_addr] <= queue_bits_wb_is_ds__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_89_en & queue_bits_wb_is_ds__T_89_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_89_addr] <= queue_bits_wb_is_ds__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_90_en & queue_bits_wb_is_ds__T_90_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_90_addr] <= queue_bits_wb_is_ds__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_91_en & queue_bits_wb_is_ds__T_91_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_91_addr] <= queue_bits_wb_is_ds__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_92_en & queue_bits_wb_is_ds__T_92_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_92_addr] <= queue_bits_wb_is_ds__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_93_en & queue_bits_wb_is_ds__T_93_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_93_addr] <= queue_bits_wb_is_ds__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_94_en & queue_bits_wb_is_ds__T_94_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_94_addr] <= queue_bits_wb_is_ds__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_95_en & queue_bits_wb_is_ds__T_95_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_95_addr] <= queue_bits_wb_is_ds__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_96_en & queue_bits_wb_is_ds__T_96_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_96_addr] <= queue_bits_wb_is_ds__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_97_en & queue_bits_wb_is_ds__T_97_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_97_addr] <= queue_bits_wb_is_ds__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_98_en & queue_bits_wb_is_ds__T_98_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_98_addr] <= queue_bits_wb_is_ds__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_99_en & queue_bits_wb_is_ds__T_99_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_99_addr] <= queue_bits_wb_is_ds__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_100_en & queue_bits_wb_is_ds__T_100_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_100_addr] <= queue_bits_wb_is_ds__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_101_en & queue_bits_wb_is_ds__T_101_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_101_addr] <= queue_bits_wb_is_ds__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_102_en & queue_bits_wb_is_ds__T_102_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_102_addr] <= queue_bits_wb_is_ds__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_103_en & queue_bits_wb_is_ds__T_103_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_103_addr] <= queue_bits_wb_is_ds__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_104_en & queue_bits_wb_is_ds__T_104_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_104_addr] <= queue_bits_wb_is_ds__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_105_en & queue_bits_wb_is_ds__T_105_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_105_addr] <= queue_bits_wb_is_ds__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_106_en & queue_bits_wb_is_ds__T_106_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_106_addr] <= queue_bits_wb_is_ds__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_107_en & queue_bits_wb_is_ds__T_107_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_107_addr] <= queue_bits_wb_is_ds__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_108_en & queue_bits_wb_is_ds__T_108_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_108_addr] <= queue_bits_wb_is_ds__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_109_en & queue_bits_wb_is_ds__T_109_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_109_addr] <= queue_bits_wb_is_ds__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_110_en & queue_bits_wb_is_ds__T_110_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_110_addr] <= queue_bits_wb_is_ds__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_111_en & queue_bits_wb_is_ds__T_111_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_111_addr] <= queue_bits_wb_is_ds__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_112_en & queue_bits_wb_is_ds__T_112_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_112_addr] <= queue_bits_wb_is_ds__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_113_en & queue_bits_wb_is_ds__T_113_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_113_addr] <= queue_bits_wb_is_ds__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_114_en & queue_bits_wb_is_ds__T_114_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_114_addr] <= queue_bits_wb_is_ds__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_115_en & queue_bits_wb_is_ds__T_115_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_115_addr] <= queue_bits_wb_is_ds__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_116_en & queue_bits_wb_is_ds__T_116_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_116_addr] <= queue_bits_wb_is_ds__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_117_en & queue_bits_wb_is_ds__T_117_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_117_addr] <= queue_bits_wb_is_ds__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_118_en & queue_bits_wb_is_ds__T_118_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_118_addr] <= queue_bits_wb_is_ds__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_119_en & queue_bits_wb_is_ds__T_119_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_119_addr] <= queue_bits_wb_is_ds__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_120_en & queue_bits_wb_is_ds__T_120_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_120_addr] <= queue_bits_wb_is_ds__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_121_en & queue_bits_wb_is_ds__T_121_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_121_addr] <= queue_bits_wb_is_ds__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_122_en & queue_bits_wb_is_ds__T_122_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_122_addr] <= queue_bits_wb_is_ds__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_123_en & queue_bits_wb_is_ds__T_123_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_123_addr] <= queue_bits_wb_is_ds__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_124_en & queue_bits_wb_is_ds__T_124_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_124_addr] <= queue_bits_wb_is_ds__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_125_en & queue_bits_wb_is_ds__T_125_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_125_addr] <= queue_bits_wb_is_ds__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_126_en & queue_bits_wb_is_ds__T_126_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_126_addr] <= queue_bits_wb_is_ds__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_127_en & queue_bits_wb_is_ds__T_127_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_127_addr] <= queue_bits_wb_is_ds__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_128_en & queue_bits_wb_is_ds__T_128_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_128_addr] <= queue_bits_wb_is_ds__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_129_en & queue_bits_wb_is_ds__T_129_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_129_addr] <= queue_bits_wb_is_ds__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_130_en & queue_bits_wb_is_ds__T_130_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_130_addr] <= queue_bits_wb_is_ds__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_131_en & queue_bits_wb_is_ds__T_131_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_131_addr] <= queue_bits_wb_is_ds__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_132_en & queue_bits_wb_is_ds__T_132_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_132_addr] <= queue_bits_wb_is_ds__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds__T_133_en & queue_bits_wb_is_ds__T_133_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds__T_133_addr] <= queue_bits_wb_is_ds__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_ds_q_head_w_en & queue_bits_wb_is_ds_q_head_w_mask) begin
      queue_bits_wb_is_ds[queue_bits_wb_is_ds_q_head_w_addr] <= queue_bits_wb_is_ds_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_3_en & queue_bits_wb_is_br__T_3_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_3_addr] <= queue_bits_wb_is_br__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_4_en & queue_bits_wb_is_br__T_4_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_4_addr] <= queue_bits_wb_is_br__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_5_en & queue_bits_wb_is_br__T_5_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_5_addr] <= queue_bits_wb_is_br__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_6_en & queue_bits_wb_is_br__T_6_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_6_addr] <= queue_bits_wb_is_br__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_7_en & queue_bits_wb_is_br__T_7_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_7_addr] <= queue_bits_wb_is_br__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_8_en & queue_bits_wb_is_br__T_8_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_8_addr] <= queue_bits_wb_is_br__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_9_en & queue_bits_wb_is_br__T_9_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_9_addr] <= queue_bits_wb_is_br__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_10_en & queue_bits_wb_is_br__T_10_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_10_addr] <= queue_bits_wb_is_br__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_11_en & queue_bits_wb_is_br__T_11_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_11_addr] <= queue_bits_wb_is_br__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_12_en & queue_bits_wb_is_br__T_12_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_12_addr] <= queue_bits_wb_is_br__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_13_en & queue_bits_wb_is_br__T_13_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_13_addr] <= queue_bits_wb_is_br__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_14_en & queue_bits_wb_is_br__T_14_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_14_addr] <= queue_bits_wb_is_br__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_15_en & queue_bits_wb_is_br__T_15_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_15_addr] <= queue_bits_wb_is_br__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_16_en & queue_bits_wb_is_br__T_16_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_16_addr] <= queue_bits_wb_is_br__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_17_en & queue_bits_wb_is_br__T_17_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_17_addr] <= queue_bits_wb_is_br__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_18_en & queue_bits_wb_is_br__T_18_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_18_addr] <= queue_bits_wb_is_br__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_19_en & queue_bits_wb_is_br__T_19_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_19_addr] <= queue_bits_wb_is_br__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_20_en & queue_bits_wb_is_br__T_20_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_20_addr] <= queue_bits_wb_is_br__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_21_en & queue_bits_wb_is_br__T_21_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_21_addr] <= queue_bits_wb_is_br__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_22_en & queue_bits_wb_is_br__T_22_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_22_addr] <= queue_bits_wb_is_br__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_23_en & queue_bits_wb_is_br__T_23_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_23_addr] <= queue_bits_wb_is_br__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_24_en & queue_bits_wb_is_br__T_24_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_24_addr] <= queue_bits_wb_is_br__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_25_en & queue_bits_wb_is_br__T_25_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_25_addr] <= queue_bits_wb_is_br__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_26_en & queue_bits_wb_is_br__T_26_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_26_addr] <= queue_bits_wb_is_br__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_27_en & queue_bits_wb_is_br__T_27_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_27_addr] <= queue_bits_wb_is_br__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_28_en & queue_bits_wb_is_br__T_28_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_28_addr] <= queue_bits_wb_is_br__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_29_en & queue_bits_wb_is_br__T_29_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_29_addr] <= queue_bits_wb_is_br__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_30_en & queue_bits_wb_is_br__T_30_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_30_addr] <= queue_bits_wb_is_br__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_31_en & queue_bits_wb_is_br__T_31_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_31_addr] <= queue_bits_wb_is_br__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_32_en & queue_bits_wb_is_br__T_32_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_32_addr] <= queue_bits_wb_is_br__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_33_en & queue_bits_wb_is_br__T_33_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_33_addr] <= queue_bits_wb_is_br__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_34_en & queue_bits_wb_is_br__T_34_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_34_addr] <= queue_bits_wb_is_br__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_35_en & queue_bits_wb_is_br__T_35_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_35_addr] <= queue_bits_wb_is_br__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_36_en & queue_bits_wb_is_br__T_36_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_36_addr] <= queue_bits_wb_is_br__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_37_en & queue_bits_wb_is_br__T_37_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_37_addr] <= queue_bits_wb_is_br__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_38_en & queue_bits_wb_is_br__T_38_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_38_addr] <= queue_bits_wb_is_br__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_39_en & queue_bits_wb_is_br__T_39_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_39_addr] <= queue_bits_wb_is_br__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_40_en & queue_bits_wb_is_br__T_40_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_40_addr] <= queue_bits_wb_is_br__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_41_en & queue_bits_wb_is_br__T_41_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_41_addr] <= queue_bits_wb_is_br__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_42_en & queue_bits_wb_is_br__T_42_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_42_addr] <= queue_bits_wb_is_br__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_43_en & queue_bits_wb_is_br__T_43_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_43_addr] <= queue_bits_wb_is_br__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_44_en & queue_bits_wb_is_br__T_44_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_44_addr] <= queue_bits_wb_is_br__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_45_en & queue_bits_wb_is_br__T_45_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_45_addr] <= queue_bits_wb_is_br__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_46_en & queue_bits_wb_is_br__T_46_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_46_addr] <= queue_bits_wb_is_br__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_47_en & queue_bits_wb_is_br__T_47_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_47_addr] <= queue_bits_wb_is_br__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_48_en & queue_bits_wb_is_br__T_48_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_48_addr] <= queue_bits_wb_is_br__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_49_en & queue_bits_wb_is_br__T_49_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_49_addr] <= queue_bits_wb_is_br__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_50_en & queue_bits_wb_is_br__T_50_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_50_addr] <= queue_bits_wb_is_br__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_51_en & queue_bits_wb_is_br__T_51_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_51_addr] <= queue_bits_wb_is_br__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_52_en & queue_bits_wb_is_br__T_52_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_52_addr] <= queue_bits_wb_is_br__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_53_en & queue_bits_wb_is_br__T_53_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_53_addr] <= queue_bits_wb_is_br__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_54_en & queue_bits_wb_is_br__T_54_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_54_addr] <= queue_bits_wb_is_br__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_55_en & queue_bits_wb_is_br__T_55_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_55_addr] <= queue_bits_wb_is_br__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_56_en & queue_bits_wb_is_br__T_56_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_56_addr] <= queue_bits_wb_is_br__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_57_en & queue_bits_wb_is_br__T_57_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_57_addr] <= queue_bits_wb_is_br__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_58_en & queue_bits_wb_is_br__T_58_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_58_addr] <= queue_bits_wb_is_br__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_59_en & queue_bits_wb_is_br__T_59_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_59_addr] <= queue_bits_wb_is_br__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_60_en & queue_bits_wb_is_br__T_60_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_60_addr] <= queue_bits_wb_is_br__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_61_en & queue_bits_wb_is_br__T_61_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_61_addr] <= queue_bits_wb_is_br__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_62_en & queue_bits_wb_is_br__T_62_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_62_addr] <= queue_bits_wb_is_br__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_63_en & queue_bits_wb_is_br__T_63_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_63_addr] <= queue_bits_wb_is_br__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_64_en & queue_bits_wb_is_br__T_64_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_64_addr] <= queue_bits_wb_is_br__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_65_en & queue_bits_wb_is_br__T_65_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_65_addr] <= queue_bits_wb_is_br__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_66_en & queue_bits_wb_is_br__T_66_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_66_addr] <= queue_bits_wb_is_br__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_67_en & queue_bits_wb_is_br__T_67_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_67_addr] <= queue_bits_wb_is_br__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_68_en & queue_bits_wb_is_br__T_68_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_68_addr] <= queue_bits_wb_is_br__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_70_en & queue_bits_wb_is_br__T_70_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_70_addr] <= queue_bits_wb_is_br__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_71_en & queue_bits_wb_is_br__T_71_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_71_addr] <= queue_bits_wb_is_br__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_72_en & queue_bits_wb_is_br__T_72_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_72_addr] <= queue_bits_wb_is_br__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_73_en & queue_bits_wb_is_br__T_73_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_73_addr] <= queue_bits_wb_is_br__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_74_en & queue_bits_wb_is_br__T_74_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_74_addr] <= queue_bits_wb_is_br__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_75_en & queue_bits_wb_is_br__T_75_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_75_addr] <= queue_bits_wb_is_br__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_76_en & queue_bits_wb_is_br__T_76_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_76_addr] <= queue_bits_wb_is_br__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_77_en & queue_bits_wb_is_br__T_77_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_77_addr] <= queue_bits_wb_is_br__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_78_en & queue_bits_wb_is_br__T_78_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_78_addr] <= queue_bits_wb_is_br__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_79_en & queue_bits_wb_is_br__T_79_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_79_addr] <= queue_bits_wb_is_br__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_80_en & queue_bits_wb_is_br__T_80_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_80_addr] <= queue_bits_wb_is_br__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_81_en & queue_bits_wb_is_br__T_81_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_81_addr] <= queue_bits_wb_is_br__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_82_en & queue_bits_wb_is_br__T_82_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_82_addr] <= queue_bits_wb_is_br__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_83_en & queue_bits_wb_is_br__T_83_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_83_addr] <= queue_bits_wb_is_br__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_84_en & queue_bits_wb_is_br__T_84_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_84_addr] <= queue_bits_wb_is_br__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_85_en & queue_bits_wb_is_br__T_85_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_85_addr] <= queue_bits_wb_is_br__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_86_en & queue_bits_wb_is_br__T_86_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_86_addr] <= queue_bits_wb_is_br__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_87_en & queue_bits_wb_is_br__T_87_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_87_addr] <= queue_bits_wb_is_br__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_88_en & queue_bits_wb_is_br__T_88_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_88_addr] <= queue_bits_wb_is_br__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_89_en & queue_bits_wb_is_br__T_89_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_89_addr] <= queue_bits_wb_is_br__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_90_en & queue_bits_wb_is_br__T_90_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_90_addr] <= queue_bits_wb_is_br__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_91_en & queue_bits_wb_is_br__T_91_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_91_addr] <= queue_bits_wb_is_br__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_92_en & queue_bits_wb_is_br__T_92_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_92_addr] <= queue_bits_wb_is_br__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_93_en & queue_bits_wb_is_br__T_93_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_93_addr] <= queue_bits_wb_is_br__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_94_en & queue_bits_wb_is_br__T_94_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_94_addr] <= queue_bits_wb_is_br__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_95_en & queue_bits_wb_is_br__T_95_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_95_addr] <= queue_bits_wb_is_br__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_96_en & queue_bits_wb_is_br__T_96_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_96_addr] <= queue_bits_wb_is_br__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_97_en & queue_bits_wb_is_br__T_97_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_97_addr] <= queue_bits_wb_is_br__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_98_en & queue_bits_wb_is_br__T_98_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_98_addr] <= queue_bits_wb_is_br__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_99_en & queue_bits_wb_is_br__T_99_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_99_addr] <= queue_bits_wb_is_br__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_100_en & queue_bits_wb_is_br__T_100_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_100_addr] <= queue_bits_wb_is_br__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_101_en & queue_bits_wb_is_br__T_101_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_101_addr] <= queue_bits_wb_is_br__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_102_en & queue_bits_wb_is_br__T_102_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_102_addr] <= queue_bits_wb_is_br__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_103_en & queue_bits_wb_is_br__T_103_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_103_addr] <= queue_bits_wb_is_br__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_104_en & queue_bits_wb_is_br__T_104_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_104_addr] <= queue_bits_wb_is_br__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_105_en & queue_bits_wb_is_br__T_105_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_105_addr] <= queue_bits_wb_is_br__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_106_en & queue_bits_wb_is_br__T_106_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_106_addr] <= queue_bits_wb_is_br__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_107_en & queue_bits_wb_is_br__T_107_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_107_addr] <= queue_bits_wb_is_br__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_108_en & queue_bits_wb_is_br__T_108_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_108_addr] <= queue_bits_wb_is_br__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_109_en & queue_bits_wb_is_br__T_109_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_109_addr] <= queue_bits_wb_is_br__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_110_en & queue_bits_wb_is_br__T_110_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_110_addr] <= queue_bits_wb_is_br__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_111_en & queue_bits_wb_is_br__T_111_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_111_addr] <= queue_bits_wb_is_br__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_112_en & queue_bits_wb_is_br__T_112_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_112_addr] <= queue_bits_wb_is_br__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_113_en & queue_bits_wb_is_br__T_113_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_113_addr] <= queue_bits_wb_is_br__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_114_en & queue_bits_wb_is_br__T_114_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_114_addr] <= queue_bits_wb_is_br__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_115_en & queue_bits_wb_is_br__T_115_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_115_addr] <= queue_bits_wb_is_br__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_116_en & queue_bits_wb_is_br__T_116_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_116_addr] <= queue_bits_wb_is_br__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_117_en & queue_bits_wb_is_br__T_117_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_117_addr] <= queue_bits_wb_is_br__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_118_en & queue_bits_wb_is_br__T_118_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_118_addr] <= queue_bits_wb_is_br__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_119_en & queue_bits_wb_is_br__T_119_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_119_addr] <= queue_bits_wb_is_br__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_120_en & queue_bits_wb_is_br__T_120_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_120_addr] <= queue_bits_wb_is_br__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_121_en & queue_bits_wb_is_br__T_121_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_121_addr] <= queue_bits_wb_is_br__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_122_en & queue_bits_wb_is_br__T_122_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_122_addr] <= queue_bits_wb_is_br__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_123_en & queue_bits_wb_is_br__T_123_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_123_addr] <= queue_bits_wb_is_br__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_124_en & queue_bits_wb_is_br__T_124_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_124_addr] <= queue_bits_wb_is_br__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_125_en & queue_bits_wb_is_br__T_125_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_125_addr] <= queue_bits_wb_is_br__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_126_en & queue_bits_wb_is_br__T_126_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_126_addr] <= queue_bits_wb_is_br__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_127_en & queue_bits_wb_is_br__T_127_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_127_addr] <= queue_bits_wb_is_br__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_128_en & queue_bits_wb_is_br__T_128_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_128_addr] <= queue_bits_wb_is_br__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_129_en & queue_bits_wb_is_br__T_129_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_129_addr] <= queue_bits_wb_is_br__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_130_en & queue_bits_wb_is_br__T_130_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_130_addr] <= queue_bits_wb_is_br__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_131_en & queue_bits_wb_is_br__T_131_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_131_addr] <= queue_bits_wb_is_br__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_132_en & queue_bits_wb_is_br__T_132_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_132_addr] <= queue_bits_wb_is_br__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br__T_133_en & queue_bits_wb_is_br__T_133_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br__T_133_addr] <= queue_bits_wb_is_br__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_is_br_q_head_w_en & queue_bits_wb_is_br_q_head_w_mask) begin
      queue_bits_wb_is_br[queue_bits_wb_is_br_q_head_w_addr] <= queue_bits_wb_is_br_q_head_w_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_3_en & queue_bits_wb_npc__T_3_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_3_addr] <= queue_bits_wb_npc__T_3_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_4_en & queue_bits_wb_npc__T_4_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_4_addr] <= queue_bits_wb_npc__T_4_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_5_en & queue_bits_wb_npc__T_5_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_5_addr] <= queue_bits_wb_npc__T_5_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_6_en & queue_bits_wb_npc__T_6_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_6_addr] <= queue_bits_wb_npc__T_6_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_7_en & queue_bits_wb_npc__T_7_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_7_addr] <= queue_bits_wb_npc__T_7_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_8_en & queue_bits_wb_npc__T_8_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_8_addr] <= queue_bits_wb_npc__T_8_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_9_en & queue_bits_wb_npc__T_9_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_9_addr] <= queue_bits_wb_npc__T_9_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_10_en & queue_bits_wb_npc__T_10_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_10_addr] <= queue_bits_wb_npc__T_10_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_11_en & queue_bits_wb_npc__T_11_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_11_addr] <= queue_bits_wb_npc__T_11_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_12_en & queue_bits_wb_npc__T_12_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_12_addr] <= queue_bits_wb_npc__T_12_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_13_en & queue_bits_wb_npc__T_13_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_13_addr] <= queue_bits_wb_npc__T_13_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_14_en & queue_bits_wb_npc__T_14_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_14_addr] <= queue_bits_wb_npc__T_14_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_15_en & queue_bits_wb_npc__T_15_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_15_addr] <= queue_bits_wb_npc__T_15_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_16_en & queue_bits_wb_npc__T_16_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_16_addr] <= queue_bits_wb_npc__T_16_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_17_en & queue_bits_wb_npc__T_17_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_17_addr] <= queue_bits_wb_npc__T_17_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_18_en & queue_bits_wb_npc__T_18_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_18_addr] <= queue_bits_wb_npc__T_18_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_19_en & queue_bits_wb_npc__T_19_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_19_addr] <= queue_bits_wb_npc__T_19_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_20_en & queue_bits_wb_npc__T_20_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_20_addr] <= queue_bits_wb_npc__T_20_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_21_en & queue_bits_wb_npc__T_21_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_21_addr] <= queue_bits_wb_npc__T_21_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_22_en & queue_bits_wb_npc__T_22_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_22_addr] <= queue_bits_wb_npc__T_22_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_23_en & queue_bits_wb_npc__T_23_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_23_addr] <= queue_bits_wb_npc__T_23_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_24_en & queue_bits_wb_npc__T_24_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_24_addr] <= queue_bits_wb_npc__T_24_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_25_en & queue_bits_wb_npc__T_25_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_25_addr] <= queue_bits_wb_npc__T_25_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_26_en & queue_bits_wb_npc__T_26_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_26_addr] <= queue_bits_wb_npc__T_26_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_27_en & queue_bits_wb_npc__T_27_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_27_addr] <= queue_bits_wb_npc__T_27_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_28_en & queue_bits_wb_npc__T_28_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_28_addr] <= queue_bits_wb_npc__T_28_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_29_en & queue_bits_wb_npc__T_29_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_29_addr] <= queue_bits_wb_npc__T_29_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_30_en & queue_bits_wb_npc__T_30_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_30_addr] <= queue_bits_wb_npc__T_30_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_31_en & queue_bits_wb_npc__T_31_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_31_addr] <= queue_bits_wb_npc__T_31_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_32_en & queue_bits_wb_npc__T_32_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_32_addr] <= queue_bits_wb_npc__T_32_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_33_en & queue_bits_wb_npc__T_33_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_33_addr] <= queue_bits_wb_npc__T_33_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_34_en & queue_bits_wb_npc__T_34_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_34_addr] <= queue_bits_wb_npc__T_34_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_35_en & queue_bits_wb_npc__T_35_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_35_addr] <= queue_bits_wb_npc__T_35_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_36_en & queue_bits_wb_npc__T_36_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_36_addr] <= queue_bits_wb_npc__T_36_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_37_en & queue_bits_wb_npc__T_37_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_37_addr] <= queue_bits_wb_npc__T_37_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_38_en & queue_bits_wb_npc__T_38_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_38_addr] <= queue_bits_wb_npc__T_38_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_39_en & queue_bits_wb_npc__T_39_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_39_addr] <= queue_bits_wb_npc__T_39_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_40_en & queue_bits_wb_npc__T_40_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_40_addr] <= queue_bits_wb_npc__T_40_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_41_en & queue_bits_wb_npc__T_41_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_41_addr] <= queue_bits_wb_npc__T_41_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_42_en & queue_bits_wb_npc__T_42_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_42_addr] <= queue_bits_wb_npc__T_42_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_43_en & queue_bits_wb_npc__T_43_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_43_addr] <= queue_bits_wb_npc__T_43_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_44_en & queue_bits_wb_npc__T_44_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_44_addr] <= queue_bits_wb_npc__T_44_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_45_en & queue_bits_wb_npc__T_45_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_45_addr] <= queue_bits_wb_npc__T_45_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_46_en & queue_bits_wb_npc__T_46_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_46_addr] <= queue_bits_wb_npc__T_46_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_47_en & queue_bits_wb_npc__T_47_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_47_addr] <= queue_bits_wb_npc__T_47_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_48_en & queue_bits_wb_npc__T_48_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_48_addr] <= queue_bits_wb_npc__T_48_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_49_en & queue_bits_wb_npc__T_49_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_49_addr] <= queue_bits_wb_npc__T_49_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_50_en & queue_bits_wb_npc__T_50_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_50_addr] <= queue_bits_wb_npc__T_50_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_51_en & queue_bits_wb_npc__T_51_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_51_addr] <= queue_bits_wb_npc__T_51_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_52_en & queue_bits_wb_npc__T_52_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_52_addr] <= queue_bits_wb_npc__T_52_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_53_en & queue_bits_wb_npc__T_53_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_53_addr] <= queue_bits_wb_npc__T_53_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_54_en & queue_bits_wb_npc__T_54_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_54_addr] <= queue_bits_wb_npc__T_54_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_55_en & queue_bits_wb_npc__T_55_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_55_addr] <= queue_bits_wb_npc__T_55_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_56_en & queue_bits_wb_npc__T_56_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_56_addr] <= queue_bits_wb_npc__T_56_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_57_en & queue_bits_wb_npc__T_57_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_57_addr] <= queue_bits_wb_npc__T_57_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_58_en & queue_bits_wb_npc__T_58_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_58_addr] <= queue_bits_wb_npc__T_58_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_59_en & queue_bits_wb_npc__T_59_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_59_addr] <= queue_bits_wb_npc__T_59_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_60_en & queue_bits_wb_npc__T_60_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_60_addr] <= queue_bits_wb_npc__T_60_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_61_en & queue_bits_wb_npc__T_61_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_61_addr] <= queue_bits_wb_npc__T_61_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_62_en & queue_bits_wb_npc__T_62_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_62_addr] <= queue_bits_wb_npc__T_62_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_63_en & queue_bits_wb_npc__T_63_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_63_addr] <= queue_bits_wb_npc__T_63_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_64_en & queue_bits_wb_npc__T_64_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_64_addr] <= queue_bits_wb_npc__T_64_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_65_en & queue_bits_wb_npc__T_65_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_65_addr] <= queue_bits_wb_npc__T_65_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_66_en & queue_bits_wb_npc__T_66_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_66_addr] <= queue_bits_wb_npc__T_66_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_67_en & queue_bits_wb_npc__T_67_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_67_addr] <= queue_bits_wb_npc__T_67_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_68_en & queue_bits_wb_npc__T_68_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_68_addr] <= queue_bits_wb_npc__T_68_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_70_en & queue_bits_wb_npc__T_70_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_70_addr] <= queue_bits_wb_npc__T_70_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_71_en & queue_bits_wb_npc__T_71_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_71_addr] <= queue_bits_wb_npc__T_71_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_72_en & queue_bits_wb_npc__T_72_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_72_addr] <= queue_bits_wb_npc__T_72_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_73_en & queue_bits_wb_npc__T_73_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_73_addr] <= queue_bits_wb_npc__T_73_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_74_en & queue_bits_wb_npc__T_74_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_74_addr] <= queue_bits_wb_npc__T_74_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_75_en & queue_bits_wb_npc__T_75_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_75_addr] <= queue_bits_wb_npc__T_75_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_76_en & queue_bits_wb_npc__T_76_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_76_addr] <= queue_bits_wb_npc__T_76_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_77_en & queue_bits_wb_npc__T_77_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_77_addr] <= queue_bits_wb_npc__T_77_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_78_en & queue_bits_wb_npc__T_78_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_78_addr] <= queue_bits_wb_npc__T_78_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_79_en & queue_bits_wb_npc__T_79_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_79_addr] <= queue_bits_wb_npc__T_79_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_80_en & queue_bits_wb_npc__T_80_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_80_addr] <= queue_bits_wb_npc__T_80_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_81_en & queue_bits_wb_npc__T_81_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_81_addr] <= queue_bits_wb_npc__T_81_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_82_en & queue_bits_wb_npc__T_82_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_82_addr] <= queue_bits_wb_npc__T_82_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_83_en & queue_bits_wb_npc__T_83_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_83_addr] <= queue_bits_wb_npc__T_83_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_84_en & queue_bits_wb_npc__T_84_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_84_addr] <= queue_bits_wb_npc__T_84_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_85_en & queue_bits_wb_npc__T_85_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_85_addr] <= queue_bits_wb_npc__T_85_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_86_en & queue_bits_wb_npc__T_86_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_86_addr] <= queue_bits_wb_npc__T_86_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_87_en & queue_bits_wb_npc__T_87_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_87_addr] <= queue_bits_wb_npc__T_87_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_88_en & queue_bits_wb_npc__T_88_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_88_addr] <= queue_bits_wb_npc__T_88_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_89_en & queue_bits_wb_npc__T_89_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_89_addr] <= queue_bits_wb_npc__T_89_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_90_en & queue_bits_wb_npc__T_90_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_90_addr] <= queue_bits_wb_npc__T_90_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_91_en & queue_bits_wb_npc__T_91_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_91_addr] <= queue_bits_wb_npc__T_91_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_92_en & queue_bits_wb_npc__T_92_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_92_addr] <= queue_bits_wb_npc__T_92_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_93_en & queue_bits_wb_npc__T_93_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_93_addr] <= queue_bits_wb_npc__T_93_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_94_en & queue_bits_wb_npc__T_94_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_94_addr] <= queue_bits_wb_npc__T_94_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_95_en & queue_bits_wb_npc__T_95_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_95_addr] <= queue_bits_wb_npc__T_95_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_96_en & queue_bits_wb_npc__T_96_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_96_addr] <= queue_bits_wb_npc__T_96_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_97_en & queue_bits_wb_npc__T_97_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_97_addr] <= queue_bits_wb_npc__T_97_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_98_en & queue_bits_wb_npc__T_98_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_98_addr] <= queue_bits_wb_npc__T_98_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_99_en & queue_bits_wb_npc__T_99_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_99_addr] <= queue_bits_wb_npc__T_99_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_100_en & queue_bits_wb_npc__T_100_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_100_addr] <= queue_bits_wb_npc__T_100_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_101_en & queue_bits_wb_npc__T_101_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_101_addr] <= queue_bits_wb_npc__T_101_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_102_en & queue_bits_wb_npc__T_102_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_102_addr] <= queue_bits_wb_npc__T_102_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_103_en & queue_bits_wb_npc__T_103_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_103_addr] <= queue_bits_wb_npc__T_103_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_104_en & queue_bits_wb_npc__T_104_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_104_addr] <= queue_bits_wb_npc__T_104_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_105_en & queue_bits_wb_npc__T_105_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_105_addr] <= queue_bits_wb_npc__T_105_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_106_en & queue_bits_wb_npc__T_106_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_106_addr] <= queue_bits_wb_npc__T_106_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_107_en & queue_bits_wb_npc__T_107_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_107_addr] <= queue_bits_wb_npc__T_107_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_108_en & queue_bits_wb_npc__T_108_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_108_addr] <= queue_bits_wb_npc__T_108_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_109_en & queue_bits_wb_npc__T_109_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_109_addr] <= queue_bits_wb_npc__T_109_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_110_en & queue_bits_wb_npc__T_110_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_110_addr] <= queue_bits_wb_npc__T_110_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_111_en & queue_bits_wb_npc__T_111_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_111_addr] <= queue_bits_wb_npc__T_111_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_112_en & queue_bits_wb_npc__T_112_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_112_addr] <= queue_bits_wb_npc__T_112_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_113_en & queue_bits_wb_npc__T_113_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_113_addr] <= queue_bits_wb_npc__T_113_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_114_en & queue_bits_wb_npc__T_114_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_114_addr] <= queue_bits_wb_npc__T_114_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_115_en & queue_bits_wb_npc__T_115_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_115_addr] <= queue_bits_wb_npc__T_115_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_116_en & queue_bits_wb_npc__T_116_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_116_addr] <= queue_bits_wb_npc__T_116_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_117_en & queue_bits_wb_npc__T_117_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_117_addr] <= queue_bits_wb_npc__T_117_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_118_en & queue_bits_wb_npc__T_118_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_118_addr] <= queue_bits_wb_npc__T_118_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_119_en & queue_bits_wb_npc__T_119_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_119_addr] <= queue_bits_wb_npc__T_119_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_120_en & queue_bits_wb_npc__T_120_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_120_addr] <= queue_bits_wb_npc__T_120_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_121_en & queue_bits_wb_npc__T_121_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_121_addr] <= queue_bits_wb_npc__T_121_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_122_en & queue_bits_wb_npc__T_122_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_122_addr] <= queue_bits_wb_npc__T_122_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_123_en & queue_bits_wb_npc__T_123_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_123_addr] <= queue_bits_wb_npc__T_123_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_124_en & queue_bits_wb_npc__T_124_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_124_addr] <= queue_bits_wb_npc__T_124_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_125_en & queue_bits_wb_npc__T_125_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_125_addr] <= queue_bits_wb_npc__T_125_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_126_en & queue_bits_wb_npc__T_126_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_126_addr] <= queue_bits_wb_npc__T_126_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_127_en & queue_bits_wb_npc__T_127_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_127_addr] <= queue_bits_wb_npc__T_127_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_128_en & queue_bits_wb_npc__T_128_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_128_addr] <= queue_bits_wb_npc__T_128_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_129_en & queue_bits_wb_npc__T_129_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_129_addr] <= queue_bits_wb_npc__T_129_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_130_en & queue_bits_wb_npc__T_130_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_130_addr] <= queue_bits_wb_npc__T_130_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_131_en & queue_bits_wb_npc__T_131_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_131_addr] <= queue_bits_wb_npc__T_131_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_132_en & queue_bits_wb_npc__T_132_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_132_addr] <= queue_bits_wb_npc__T_132_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc__T_133_en & queue_bits_wb_npc__T_133_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc__T_133_addr] <= queue_bits_wb_npc__T_133_data; // @[utils.scala 30:18]
    end
    if(queue_bits_wb_npc_q_head_w_en & queue_bits_wb_npc_q_head_w_mask) begin
      queue_bits_wb_npc[queue_bits_wb_npc_q_head_w_addr] <= queue_bits_wb_npc_q_head_w_data; // @[utils.scala 30:18]
    end
    if (reset) begin
      head <= 6'h0;
    end else if (io_deq_valid) begin
      head <= _T_2;
    end
  end
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_ip7,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  input  [4:0]  io_fu_in_bits_ops_fu_op,
  input  [31:0] io_fu_in_bits_ops_op1,
  input  [31:0] io_fu_in_bits_ops_op2,
  output        io_fu_out_valid,
  output        io_fu_out_bits_v,
  output [7:0]  io_fu_out_bits_id,
  output [31:0] io_fu_out_bits_pc,
  output [5:0]  io_fu_out_bits_instr_op,
  output [4:0]  io_fu_out_bits_instr_rs_idx,
  output [4:0]  io_fu_out_bits_instr_rt_idx,
  output [4:0]  io_fu_out_bits_instr_rd_idx,
  output [4:0]  io_fu_out_bits_instr_shamt,
  output [5:0]  io_fu_out_bits_instr_func,
  output [4:0]  io_fu_out_bits_rd_idx,
  output        io_fu_out_bits_wen,
  output [31:0] io_fu_out_bits_data,
  output        io_fu_out_bits_ip7,
  output        io_fu_out_bits_is_ds,
  output        io_fu_out_bits_is_br,
  output [31:0] io_fu_out_bits_npc,
  output        io_working,
  output        io_divider_data_dividend_tvalid,
  output        io_divider_data_divisor_tvalid,
  input         io_divider_data_dout_tvalid,
  output [39:0] io_divider_data_dividend_tdata,
  output [39:0] io_divider_data_divisor_tdata,
  input  [79:0] io_divider_data_dout_tdata,
  output [32:0] io_multiplier_data_a,
  output [32:0] io_multiplier_data_b,
  input  [65:0] io_multiplier_data_dout
);
  wire  multiplier_clock; // @[mdu.scala 150:26]
  wire  multiplier_reset; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_in_ready; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_in_valid; // @[mdu.scala 150:26]
  wire [5:0] multiplier_io_fu_in_bits_id; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_in_bits_fu_op; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_in_bits_op1; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_in_bits_op2; // @[mdu.scala 150:26]
  wire [7:0] multiplier_io_fu_in_bits_wb_id; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_in_bits_wb_pc; // @[mdu.scala 150:26]
  wire [5:0] multiplier_io_fu_in_bits_wb_instr_op; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_in_bits_wb_instr_rs_idx; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_in_bits_wb_instr_rt_idx; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_in_bits_wb_instr_rd_idx; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_in_bits_wb_instr_shamt; // @[mdu.scala 150:26]
  wire [5:0] multiplier_io_fu_in_bits_wb_instr_func; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_in_bits_wb_rd_idx; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_in_bits_wb_ip7; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_in_bits_wb_is_ds; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_in_bits_wb_is_br; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_in_bits_wb_npc; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_out_valid; // @[mdu.scala 150:26]
  wire [5:0] multiplier_io_fu_out_bits_id; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_out_bits_hi; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_out_bits_lo; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_out_bits_op1; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_out_bits_fu_op; // @[mdu.scala 150:26]
  wire [7:0] multiplier_io_fu_out_bits_wb_id; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_out_bits_wb_pc; // @[mdu.scala 150:26]
  wire [5:0] multiplier_io_fu_out_bits_wb_instr_op; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_out_bits_wb_instr_rs_idx; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_out_bits_wb_instr_rt_idx; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_out_bits_wb_instr_rd_idx; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_out_bits_wb_instr_shamt; // @[mdu.scala 150:26]
  wire [5:0] multiplier_io_fu_out_bits_wb_instr_func; // @[mdu.scala 150:26]
  wire [4:0] multiplier_io_fu_out_bits_wb_rd_idx; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_out_bits_wb_ip7; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_out_bits_wb_is_ds; // @[mdu.scala 150:26]
  wire  multiplier_io_fu_out_bits_wb_is_br; // @[mdu.scala 150:26]
  wire [31:0] multiplier_io_fu_out_bits_wb_npc; // @[mdu.scala 150:26]
  wire [32:0] multiplier_io_multiplier_data_a; // @[mdu.scala 150:26]
  wire [32:0] multiplier_io_multiplier_data_b; // @[mdu.scala 150:26]
  wire [65:0] multiplier_io_multiplier_data_dout; // @[mdu.scala 150:26]
  wire  divider_clock; // @[mdu.scala 151:23]
  wire  divider_reset; // @[mdu.scala 151:23]
  wire  divider_io_fu_in_valid; // @[mdu.scala 151:23]
  wire [5:0] divider_io_fu_in_bits_id; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_in_bits_fu_op; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_in_bits_op1; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_in_bits_op2; // @[mdu.scala 151:23]
  wire [7:0] divider_io_fu_in_bits_wb_id; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_in_bits_wb_pc; // @[mdu.scala 151:23]
  wire [5:0] divider_io_fu_in_bits_wb_instr_op; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_in_bits_wb_instr_rs_idx; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_in_bits_wb_instr_rt_idx; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_in_bits_wb_instr_rd_idx; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_in_bits_wb_instr_shamt; // @[mdu.scala 151:23]
  wire [5:0] divider_io_fu_in_bits_wb_instr_func; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_in_bits_wb_rd_idx; // @[mdu.scala 151:23]
  wire  divider_io_fu_in_bits_wb_ip7; // @[mdu.scala 151:23]
  wire  divider_io_fu_in_bits_wb_is_ds; // @[mdu.scala 151:23]
  wire  divider_io_fu_in_bits_wb_is_br; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_in_bits_wb_npc; // @[mdu.scala 151:23]
  wire  divider_io_fu_out_valid; // @[mdu.scala 151:23]
  wire [5:0] divider_io_fu_out_bits_id; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_out_bits_hi; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_out_bits_lo; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_out_bits_op1; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_out_bits_fu_op; // @[mdu.scala 151:23]
  wire [7:0] divider_io_fu_out_bits_wb_id; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_out_bits_wb_pc; // @[mdu.scala 151:23]
  wire [5:0] divider_io_fu_out_bits_wb_instr_op; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_out_bits_wb_instr_rs_idx; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_out_bits_wb_instr_rt_idx; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_out_bits_wb_instr_rd_idx; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_out_bits_wb_instr_shamt; // @[mdu.scala 151:23]
  wire [5:0] divider_io_fu_out_bits_wb_instr_func; // @[mdu.scala 151:23]
  wire [4:0] divider_io_fu_out_bits_wb_rd_idx; // @[mdu.scala 151:23]
  wire  divider_io_fu_out_bits_wb_ip7; // @[mdu.scala 151:23]
  wire  divider_io_fu_out_bits_wb_is_ds; // @[mdu.scala 151:23]
  wire  divider_io_fu_out_bits_wb_is_br; // @[mdu.scala 151:23]
  wire [31:0] divider_io_fu_out_bits_wb_npc; // @[mdu.scala 151:23]
  wire  divider_io_divider_data_dividend_tvalid; // @[mdu.scala 151:23]
  wire  divider_io_divider_data_divisor_tvalid; // @[mdu.scala 151:23]
  wire  divider_io_divider_data_dout_tvalid; // @[mdu.scala 151:23]
  wire [39:0] divider_io_divider_data_dividend_tdata; // @[mdu.scala 151:23]
  wire [39:0] divider_io_divider_data_divisor_tdata; // @[mdu.scala 151:23]
  wire [79:0] divider_io_divider_data_dout_tdata; // @[mdu.scala 151:23]
  wire  rob_clock; // @[mdu.scala 152:19]
  wire  rob_reset; // @[mdu.scala 152:19]
  wire  rob_io_enq_0_valid; // @[mdu.scala 152:19]
  wire [5:0] rob_io_enq_0_bits_id; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_0_bits_data_hi; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_0_bits_data_lo; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_0_bits_data_op1; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_0_bits_data_fu_op; // @[mdu.scala 152:19]
  wire [7:0] rob_io_enq_0_bits_data_wb_id; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_0_bits_data_wb_pc; // @[mdu.scala 152:19]
  wire [5:0] rob_io_enq_0_bits_data_wb_instr_op; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_0_bits_data_wb_instr_rs_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_0_bits_data_wb_instr_rt_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_0_bits_data_wb_instr_rd_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_0_bits_data_wb_instr_shamt; // @[mdu.scala 152:19]
  wire [5:0] rob_io_enq_0_bits_data_wb_instr_func; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_0_bits_data_wb_rd_idx; // @[mdu.scala 152:19]
  wire  rob_io_enq_0_bits_data_wb_ip7; // @[mdu.scala 152:19]
  wire  rob_io_enq_0_bits_data_wb_is_ds; // @[mdu.scala 152:19]
  wire  rob_io_enq_0_bits_data_wb_is_br; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_0_bits_data_wb_npc; // @[mdu.scala 152:19]
  wire  rob_io_enq_1_valid; // @[mdu.scala 152:19]
  wire [5:0] rob_io_enq_1_bits_id; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_1_bits_data_hi; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_1_bits_data_lo; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_1_bits_data_op1; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_1_bits_data_fu_op; // @[mdu.scala 152:19]
  wire [7:0] rob_io_enq_1_bits_data_wb_id; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_1_bits_data_wb_pc; // @[mdu.scala 152:19]
  wire [5:0] rob_io_enq_1_bits_data_wb_instr_op; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_1_bits_data_wb_instr_rs_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_1_bits_data_wb_instr_rt_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_1_bits_data_wb_instr_rd_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_1_bits_data_wb_instr_shamt; // @[mdu.scala 152:19]
  wire [5:0] rob_io_enq_1_bits_data_wb_instr_func; // @[mdu.scala 152:19]
  wire [4:0] rob_io_enq_1_bits_data_wb_rd_idx; // @[mdu.scala 152:19]
  wire  rob_io_enq_1_bits_data_wb_ip7; // @[mdu.scala 152:19]
  wire  rob_io_enq_1_bits_data_wb_is_ds; // @[mdu.scala 152:19]
  wire  rob_io_enq_1_bits_data_wb_is_br; // @[mdu.scala 152:19]
  wire [31:0] rob_io_enq_1_bits_data_wb_npc; // @[mdu.scala 152:19]
  wire  rob_io_deq_valid; // @[mdu.scala 152:19]
  wire [31:0] rob_io_deq_bits_hi; // @[mdu.scala 152:19]
  wire [31:0] rob_io_deq_bits_lo; // @[mdu.scala 152:19]
  wire [31:0] rob_io_deq_bits_op1; // @[mdu.scala 152:19]
  wire [4:0] rob_io_deq_bits_fu_op; // @[mdu.scala 152:19]
  wire [7:0] rob_io_deq_bits_wb_id; // @[mdu.scala 152:19]
  wire [31:0] rob_io_deq_bits_wb_pc; // @[mdu.scala 152:19]
  wire [5:0] rob_io_deq_bits_wb_instr_op; // @[mdu.scala 152:19]
  wire [4:0] rob_io_deq_bits_wb_instr_rs_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_deq_bits_wb_instr_rt_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_deq_bits_wb_instr_rd_idx; // @[mdu.scala 152:19]
  wire [4:0] rob_io_deq_bits_wb_instr_shamt; // @[mdu.scala 152:19]
  wire [5:0] rob_io_deq_bits_wb_instr_func; // @[mdu.scala 152:19]
  wire [4:0] rob_io_deq_bits_wb_rd_idx; // @[mdu.scala 152:19]
  wire  rob_io_deq_bits_wb_ip7; // @[mdu.scala 152:19]
  wire  rob_io_deq_bits_wb_is_ds; // @[mdu.scala 152:19]
  wire  rob_io_deq_bits_wb_is_br; // @[mdu.scala 152:19]
  wire [31:0] rob_io_deq_bits_wb_npc; // @[mdu.scala 152:19]
  wire  _T = io_fu_in_bits_ops_fu_op == 5'hf; // @[mdu.scala 142:40]
  wire  _T_1 = io_fu_in_bits_ops_fu_op == 5'h11; // @[mdu.scala 143:29]
  wire  is_div = _T | _T_1; // @[mdu.scala 142:52]
  reg [31:0] fu_sz; // @[mdu.scala 145:22]
  reg [31:0] _RAND_0;
  reg [31:0] hi; // @[mdu.scala 147:19]
  reg [31:0] _RAND_1;
  reg [31:0] lo; // @[mdu.scala 148:19]
  reg [31:0] _RAND_2;
  reg [5:0] mduid; // @[mdu.scala 149:22]
  reg [31:0] _RAND_3;
  wire  _T_2 = ~is_div; // @[mdu.scala 155:50]
  wire  _T_7 = io_fu_in_ready & io_fu_in_valid; // @[Decoupled.scala 40:37]
  wire [5:0] _T_9 = mduid + 6'h1; // @[mdu.scala 184:43]
  wire [31:0] _GEN_3 = {{31'd0}, _T_7}; // @[mdu.scala 185:18]
  wire [31:0] _T_12 = fu_sz + _GEN_3; // @[mdu.scala 185:18]
  wire [31:0] _GEN_4 = {{31'd0}, io_fu_out_valid}; // @[mdu.scala 185:36]
  wire [31:0] _T_14 = _T_12 - _GEN_4; // @[mdu.scala 185:36]
  wire [4:0] _T_16 = rob_io_deq_bits_fu_op;
  wire  wb_rd = ~_T_16[0]; // @[mdu.scala 188:48]
  wire  wb_hilo = ~wb_rd; // @[mdu.scala 189:17]
  wire [63:0] mul = {rob_io_deq_bits_hi,rob_io_deq_bits_lo}; // @[Cat.scala 29:58]
  wire [63:0] hilo = {hi,lo}; // @[Cat.scala 29:58]
  wire  _T_19 = rob_io_deq_bits_fu_op == 5'h0; // @[mdu.scala 195:12]
  wire  _T_20 = rob_io_deq_bits_fu_op == 5'h2; // @[mdu.scala 196:12]
  wire  _T_21 = rob_io_deq_bits_fu_op == 5'h8; // @[mdu.scala 197:12]
  wire [31:0] _T_23 = _T_19 ? hi : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_24 = _T_20 ? lo : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_25 = _T_21 ? mul[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_26 = _T_23 | _T_24; // @[Mux.scala 27:72]
  wire  _T_28 = rob_io_deq_valid & wb_hilo; // @[mdu.scala 199:26]
  wire [63:0] _T_30 = hilo + mul; // @[mdu.scala 207:26]
  wire [63:0] _T_36 = hilo - mul; // @[mdu.scala 209:26]
  wire  _T_41 = 5'h19 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_43 = 5'h17 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_45 = 5'h15 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_47 = 5'h13 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_49 = 5'h11 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_51 = 5'hf == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_53 = 5'hd == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_55 = 5'hb == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_57 = 5'h7 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  wire  _T_59 = 5'h5 == rob_io_deq_bits_fu_op; // @[Mux.scala 68:19]
  MDU_Multiplier multiplier ( // @[mdu.scala 150:26]
    .clock(multiplier_clock),
    .reset(multiplier_reset),
    .io_fu_in_ready(multiplier_io_fu_in_ready),
    .io_fu_in_valid(multiplier_io_fu_in_valid),
    .io_fu_in_bits_id(multiplier_io_fu_in_bits_id),
    .io_fu_in_bits_fu_op(multiplier_io_fu_in_bits_fu_op),
    .io_fu_in_bits_op1(multiplier_io_fu_in_bits_op1),
    .io_fu_in_bits_op2(multiplier_io_fu_in_bits_op2),
    .io_fu_in_bits_wb_id(multiplier_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(multiplier_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(multiplier_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(multiplier_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(multiplier_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(multiplier_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(multiplier_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(multiplier_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(multiplier_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_ip7(multiplier_io_fu_in_bits_wb_ip7),
    .io_fu_in_bits_wb_is_ds(multiplier_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(multiplier_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(multiplier_io_fu_in_bits_wb_npc),
    .io_fu_out_valid(multiplier_io_fu_out_valid),
    .io_fu_out_bits_id(multiplier_io_fu_out_bits_id),
    .io_fu_out_bits_hi(multiplier_io_fu_out_bits_hi),
    .io_fu_out_bits_lo(multiplier_io_fu_out_bits_lo),
    .io_fu_out_bits_op1(multiplier_io_fu_out_bits_op1),
    .io_fu_out_bits_fu_op(multiplier_io_fu_out_bits_fu_op),
    .io_fu_out_bits_wb_id(multiplier_io_fu_out_bits_wb_id),
    .io_fu_out_bits_wb_pc(multiplier_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(multiplier_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(multiplier_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(multiplier_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(multiplier_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(multiplier_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(multiplier_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_rd_idx(multiplier_io_fu_out_bits_wb_rd_idx),
    .io_fu_out_bits_wb_ip7(multiplier_io_fu_out_bits_wb_ip7),
    .io_fu_out_bits_wb_is_ds(multiplier_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_wb_is_br(multiplier_io_fu_out_bits_wb_is_br),
    .io_fu_out_bits_wb_npc(multiplier_io_fu_out_bits_wb_npc),
    .io_multiplier_data_a(multiplier_io_multiplier_data_a),
    .io_multiplier_data_b(multiplier_io_multiplier_data_b),
    .io_multiplier_data_dout(multiplier_io_multiplier_data_dout)
  );
  MDU_Divider divider ( // @[mdu.scala 151:23]
    .clock(divider_clock),
    .reset(divider_reset),
    .io_fu_in_valid(divider_io_fu_in_valid),
    .io_fu_in_bits_id(divider_io_fu_in_bits_id),
    .io_fu_in_bits_fu_op(divider_io_fu_in_bits_fu_op),
    .io_fu_in_bits_op1(divider_io_fu_in_bits_op1),
    .io_fu_in_bits_op2(divider_io_fu_in_bits_op2),
    .io_fu_in_bits_wb_id(divider_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(divider_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(divider_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(divider_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(divider_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(divider_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(divider_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(divider_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(divider_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_ip7(divider_io_fu_in_bits_wb_ip7),
    .io_fu_in_bits_wb_is_ds(divider_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(divider_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(divider_io_fu_in_bits_wb_npc),
    .io_fu_out_valid(divider_io_fu_out_valid),
    .io_fu_out_bits_id(divider_io_fu_out_bits_id),
    .io_fu_out_bits_hi(divider_io_fu_out_bits_hi),
    .io_fu_out_bits_lo(divider_io_fu_out_bits_lo),
    .io_fu_out_bits_op1(divider_io_fu_out_bits_op1),
    .io_fu_out_bits_fu_op(divider_io_fu_out_bits_fu_op),
    .io_fu_out_bits_wb_id(divider_io_fu_out_bits_wb_id),
    .io_fu_out_bits_wb_pc(divider_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(divider_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(divider_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(divider_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(divider_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(divider_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(divider_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_rd_idx(divider_io_fu_out_bits_wb_rd_idx),
    .io_fu_out_bits_wb_ip7(divider_io_fu_out_bits_wb_ip7),
    .io_fu_out_bits_wb_is_ds(divider_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_wb_is_br(divider_io_fu_out_bits_wb_is_br),
    .io_fu_out_bits_wb_npc(divider_io_fu_out_bits_wb_npc),
    .io_divider_data_dividend_tvalid(divider_io_divider_data_dividend_tvalid),
    .io_divider_data_divisor_tvalid(divider_io_divider_data_divisor_tvalid),
    .io_divider_data_dout_tvalid(divider_io_divider_data_dout_tvalid),
    .io_divider_data_dividend_tdata(divider_io_divider_data_dividend_tdata),
    .io_divider_data_divisor_tdata(divider_io_divider_data_divisor_tdata),
    .io_divider_data_dout_tdata(divider_io_divider_data_dout_tdata)
  );
  ROB rob ( // @[mdu.scala 152:19]
    .clock(rob_clock),
    .reset(rob_reset),
    .io_enq_0_valid(rob_io_enq_0_valid),
    .io_enq_0_bits_id(rob_io_enq_0_bits_id),
    .io_enq_0_bits_data_hi(rob_io_enq_0_bits_data_hi),
    .io_enq_0_bits_data_lo(rob_io_enq_0_bits_data_lo),
    .io_enq_0_bits_data_op1(rob_io_enq_0_bits_data_op1),
    .io_enq_0_bits_data_fu_op(rob_io_enq_0_bits_data_fu_op),
    .io_enq_0_bits_data_wb_id(rob_io_enq_0_bits_data_wb_id),
    .io_enq_0_bits_data_wb_pc(rob_io_enq_0_bits_data_wb_pc),
    .io_enq_0_bits_data_wb_instr_op(rob_io_enq_0_bits_data_wb_instr_op),
    .io_enq_0_bits_data_wb_instr_rs_idx(rob_io_enq_0_bits_data_wb_instr_rs_idx),
    .io_enq_0_bits_data_wb_instr_rt_idx(rob_io_enq_0_bits_data_wb_instr_rt_idx),
    .io_enq_0_bits_data_wb_instr_rd_idx(rob_io_enq_0_bits_data_wb_instr_rd_idx),
    .io_enq_0_bits_data_wb_instr_shamt(rob_io_enq_0_bits_data_wb_instr_shamt),
    .io_enq_0_bits_data_wb_instr_func(rob_io_enq_0_bits_data_wb_instr_func),
    .io_enq_0_bits_data_wb_rd_idx(rob_io_enq_0_bits_data_wb_rd_idx),
    .io_enq_0_bits_data_wb_ip7(rob_io_enq_0_bits_data_wb_ip7),
    .io_enq_0_bits_data_wb_is_ds(rob_io_enq_0_bits_data_wb_is_ds),
    .io_enq_0_bits_data_wb_is_br(rob_io_enq_0_bits_data_wb_is_br),
    .io_enq_0_bits_data_wb_npc(rob_io_enq_0_bits_data_wb_npc),
    .io_enq_1_valid(rob_io_enq_1_valid),
    .io_enq_1_bits_id(rob_io_enq_1_bits_id),
    .io_enq_1_bits_data_hi(rob_io_enq_1_bits_data_hi),
    .io_enq_1_bits_data_lo(rob_io_enq_1_bits_data_lo),
    .io_enq_1_bits_data_op1(rob_io_enq_1_bits_data_op1),
    .io_enq_1_bits_data_fu_op(rob_io_enq_1_bits_data_fu_op),
    .io_enq_1_bits_data_wb_id(rob_io_enq_1_bits_data_wb_id),
    .io_enq_1_bits_data_wb_pc(rob_io_enq_1_bits_data_wb_pc),
    .io_enq_1_bits_data_wb_instr_op(rob_io_enq_1_bits_data_wb_instr_op),
    .io_enq_1_bits_data_wb_instr_rs_idx(rob_io_enq_1_bits_data_wb_instr_rs_idx),
    .io_enq_1_bits_data_wb_instr_rt_idx(rob_io_enq_1_bits_data_wb_instr_rt_idx),
    .io_enq_1_bits_data_wb_instr_rd_idx(rob_io_enq_1_bits_data_wb_instr_rd_idx),
    .io_enq_1_bits_data_wb_instr_shamt(rob_io_enq_1_bits_data_wb_instr_shamt),
    .io_enq_1_bits_data_wb_instr_func(rob_io_enq_1_bits_data_wb_instr_func),
    .io_enq_1_bits_data_wb_rd_idx(rob_io_enq_1_bits_data_wb_rd_idx),
    .io_enq_1_bits_data_wb_ip7(rob_io_enq_1_bits_data_wb_ip7),
    .io_enq_1_bits_data_wb_is_ds(rob_io_enq_1_bits_data_wb_is_ds),
    .io_enq_1_bits_data_wb_is_br(rob_io_enq_1_bits_data_wb_is_br),
    .io_enq_1_bits_data_wb_npc(rob_io_enq_1_bits_data_wb_npc),
    .io_deq_valid(rob_io_deq_valid),
    .io_deq_bits_hi(rob_io_deq_bits_hi),
    .io_deq_bits_lo(rob_io_deq_bits_lo),
    .io_deq_bits_op1(rob_io_deq_bits_op1),
    .io_deq_bits_fu_op(rob_io_deq_bits_fu_op),
    .io_deq_bits_wb_id(rob_io_deq_bits_wb_id),
    .io_deq_bits_wb_pc(rob_io_deq_bits_wb_pc),
    .io_deq_bits_wb_instr_op(rob_io_deq_bits_wb_instr_op),
    .io_deq_bits_wb_instr_rs_idx(rob_io_deq_bits_wb_instr_rs_idx),
    .io_deq_bits_wb_instr_rt_idx(rob_io_deq_bits_wb_instr_rt_idx),
    .io_deq_bits_wb_instr_rd_idx(rob_io_deq_bits_wb_instr_rd_idx),
    .io_deq_bits_wb_instr_shamt(rob_io_deq_bits_wb_instr_shamt),
    .io_deq_bits_wb_instr_func(rob_io_deq_bits_wb_instr_func),
    .io_deq_bits_wb_rd_idx(rob_io_deq_bits_wb_rd_idx),
    .io_deq_bits_wb_ip7(rob_io_deq_bits_wb_ip7),
    .io_deq_bits_wb_is_ds(rob_io_deq_bits_wb_is_ds),
    .io_deq_bits_wb_is_br(rob_io_deq_bits_wb_is_br),
    .io_deq_bits_wb_npc(rob_io_deq_bits_wb_npc)
  );
  assign io_fu_in_ready = 1'h1; // @[mdu.scala 183:18]
  assign io_fu_out_valid = rob_io_deq_valid; // @[mdu.scala 226:19]
  assign io_fu_out_bits_v = ~_T_16[0]; // @[mdu.scala 227:18 mdu.scala 228:21]
  assign io_fu_out_bits_id = rob_io_deq_bits_wb_id; // @[mdu.scala 227:18]
  assign io_fu_out_bits_pc = rob_io_deq_bits_wb_pc; // @[mdu.scala 227:18]
  assign io_fu_out_bits_instr_op = rob_io_deq_bits_wb_instr_op; // @[mdu.scala 227:18]
  assign io_fu_out_bits_instr_rs_idx = rob_io_deq_bits_wb_instr_rs_idx; // @[mdu.scala 227:18]
  assign io_fu_out_bits_instr_rt_idx = rob_io_deq_bits_wb_instr_rt_idx; // @[mdu.scala 227:18]
  assign io_fu_out_bits_instr_rd_idx = rob_io_deq_bits_wb_instr_rd_idx; // @[mdu.scala 227:18]
  assign io_fu_out_bits_instr_shamt = rob_io_deq_bits_wb_instr_shamt; // @[mdu.scala 227:18]
  assign io_fu_out_bits_instr_func = rob_io_deq_bits_wb_instr_func; // @[mdu.scala 227:18]
  assign io_fu_out_bits_rd_idx = rob_io_deq_bits_wb_rd_idx; // @[mdu.scala 227:18]
  assign io_fu_out_bits_wen = ~_T_16[0]; // @[mdu.scala 227:18 mdu.scala 229:22]
  assign io_fu_out_bits_data = _T_26 | _T_25; // @[mdu.scala 227:18 mdu.scala 230:23]
  assign io_fu_out_bits_ip7 = rob_io_deq_bits_wb_ip7; // @[mdu.scala 227:18]
  assign io_fu_out_bits_is_ds = rob_io_deq_bits_wb_is_ds; // @[mdu.scala 227:18]
  assign io_fu_out_bits_is_br = rob_io_deq_bits_wb_is_br; // @[mdu.scala 227:18]
  assign io_fu_out_bits_npc = rob_io_deq_bits_wb_npc; // @[mdu.scala 227:18]
  assign io_working = fu_sz != 32'h0; // @[mdu.scala 224:14]
  assign io_divider_data_dividend_tvalid = divider_io_divider_data_dividend_tvalid; // @[mdu.scala 170:22]
  assign io_divider_data_divisor_tvalid = divider_io_divider_data_divisor_tvalid; // @[mdu.scala 170:22]
  assign io_divider_data_dividend_tdata = divider_io_divider_data_dividend_tdata; // @[mdu.scala 170:22]
  assign io_divider_data_divisor_tdata = divider_io_divider_data_divisor_tdata; // @[mdu.scala 170:22]
  assign io_multiplier_data_a = multiplier_io_multiplier_data_a; // @[mdu.scala 161:28]
  assign io_multiplier_data_b = multiplier_io_multiplier_data_b; // @[mdu.scala 161:28]
  assign multiplier_clock = clock;
  assign multiplier_reset = reset;
  assign multiplier_io_fu_in_valid = io_fu_in_valid & _T_2; // @[mdu.scala 155:29]
  assign multiplier_io_fu_in_bits_id = mduid; // @[mdu.scala 157:31]
  assign multiplier_io_fu_in_bits_fu_op = io_fu_in_bits_ops_fu_op; // @[mdu.scala 156:34]
  assign multiplier_io_fu_in_bits_op1 = io_fu_in_bits_ops_op1; // @[mdu.scala 158:32]
  assign multiplier_io_fu_in_bits_op2 = io_fu_in_bits_ops_op2; // @[mdu.scala 159:32]
  assign multiplier_io_fu_in_bits_wb_id = io_fu_in_bits_wb_id; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_pc = io_fu_in_bits_wb_pc; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_is_ds = io_fu_in_bits_wb_is_ds; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[mdu.scala 160:31]
  assign multiplier_io_fu_in_bits_wb_npc = io_fu_in_bits_wb_npc; // @[mdu.scala 160:31]
  assign multiplier_io_multiplier_data_dout = io_multiplier_data_dout; // @[mdu.scala 161:28]
  assign divider_clock = clock;
  assign divider_reset = reset;
  assign divider_io_fu_in_valid = io_fu_in_valid & is_div; // @[mdu.scala 164:26]
  assign divider_io_fu_in_bits_id = mduid; // @[mdu.scala 166:28]
  assign divider_io_fu_in_bits_fu_op = io_fu_in_bits_ops_fu_op; // @[mdu.scala 165:31]
  assign divider_io_fu_in_bits_op1 = io_fu_in_bits_ops_op1; // @[mdu.scala 167:29]
  assign divider_io_fu_in_bits_op2 = io_fu_in_bits_ops_op2; // @[mdu.scala 168:29]
  assign divider_io_fu_in_bits_wb_id = io_fu_in_bits_wb_id; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_pc = io_fu_in_bits_wb_pc; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_is_ds = io_fu_in_bits_wb_is_ds; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[mdu.scala 169:28]
  assign divider_io_fu_in_bits_wb_npc = io_fu_in_bits_wb_npc; // @[mdu.scala 169:28]
  assign divider_io_divider_data_dout_tvalid = io_divider_data_dout_tvalid; // @[mdu.scala 170:22]
  assign divider_io_divider_data_dout_tdata = io_divider_data_dout_tdata; // @[mdu.scala 170:22]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_io_enq_0_valid = multiplier_io_fu_out_valid; // @[mdu.scala 175:23]
  assign rob_io_enq_0_bits_id = multiplier_io_fu_out_bits_id; // @[mdu.scala 176:25]
  assign rob_io_enq_0_bits_data_hi = multiplier_io_fu_out_bits_hi; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_lo = multiplier_io_fu_out_bits_lo; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_op1 = multiplier_io_fu_out_bits_op1; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_fu_op = multiplier_io_fu_out_bits_fu_op; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_id = multiplier_io_fu_out_bits_wb_id; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_pc = multiplier_io_fu_out_bits_wb_pc; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_instr_op = multiplier_io_fu_out_bits_wb_instr_op; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_instr_rs_idx = multiplier_io_fu_out_bits_wb_instr_rs_idx; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_instr_rt_idx = multiplier_io_fu_out_bits_wb_instr_rt_idx; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_instr_rd_idx = multiplier_io_fu_out_bits_wb_instr_rd_idx; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_instr_shamt = multiplier_io_fu_out_bits_wb_instr_shamt; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_instr_func = multiplier_io_fu_out_bits_wb_instr_func; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_rd_idx = multiplier_io_fu_out_bits_wb_rd_idx; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_ip7 = multiplier_io_fu_out_bits_wb_ip7; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_is_ds = multiplier_io_fu_out_bits_wb_is_ds; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_is_br = multiplier_io_fu_out_bits_wb_is_br; // @[mdu.scala 177:27]
  assign rob_io_enq_0_bits_data_wb_npc = multiplier_io_fu_out_bits_wb_npc; // @[mdu.scala 177:27]
  assign rob_io_enq_1_valid = divider_io_fu_out_valid; // @[mdu.scala 179:23]
  assign rob_io_enq_1_bits_id = divider_io_fu_out_bits_id; // @[mdu.scala 180:25]
  assign rob_io_enq_1_bits_data_hi = divider_io_fu_out_bits_hi; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_lo = divider_io_fu_out_bits_lo; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_op1 = divider_io_fu_out_bits_op1; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_fu_op = divider_io_fu_out_bits_fu_op; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_id = divider_io_fu_out_bits_wb_id; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_pc = divider_io_fu_out_bits_wb_pc; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_instr_op = divider_io_fu_out_bits_wb_instr_op; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_instr_rs_idx = divider_io_fu_out_bits_wb_instr_rs_idx; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_instr_rt_idx = divider_io_fu_out_bits_wb_instr_rt_idx; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_instr_rd_idx = divider_io_fu_out_bits_wb_instr_rd_idx; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_instr_shamt = divider_io_fu_out_bits_wb_instr_shamt; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_instr_func = divider_io_fu_out_bits_wb_instr_func; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_rd_idx = divider_io_fu_out_bits_wb_rd_idx; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_ip7 = divider_io_fu_out_bits_wb_ip7; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_is_ds = divider_io_fu_out_bits_wb_is_ds; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_is_br = divider_io_fu_out_bits_wb_is_br; // @[mdu.scala 181:27]
  assign rob_io_enq_1_bits_data_wb_npc = divider_io_fu_out_bits_wb_npc; // @[mdu.scala 181:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fu_sz = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  hi = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  lo = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mduid = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fu_sz <= 32'h0;
    end else begin
      fu_sz <= _T_14;
    end
    if (reset) begin
      hi <= 32'h0;
    end else if (_T_28) begin
      if (_T_59) begin
        hi <= rob_io_deq_bits_op1;
      end else if (!(_T_57)) begin
        if (_T_55) begin
          hi <= rob_io_deq_bits_hi;
        end else if (_T_53) begin
          hi <= rob_io_deq_bits_hi;
        end else if (_T_51) begin
          hi <= rob_io_deq_bits_hi;
        end else if (_T_49) begin
          hi <= rob_io_deq_bits_hi;
        end else if (_T_47) begin
          hi <= _T_30[63:32];
        end else if (_T_45) begin
          hi <= _T_30[63:32];
        end else if (_T_43) begin
          hi <= _T_36[63:32];
        end else if (_T_41) begin
          hi <= _T_36[63:32];
        end else begin
          hi <= 32'h0;
        end
      end
    end
    if (reset) begin
      lo <= 32'h0;
    end else if (_T_28) begin
      if (!(_T_59)) begin
        if (_T_57) begin
          lo <= rob_io_deq_bits_op1;
        end else if (_T_55) begin
          lo <= rob_io_deq_bits_lo;
        end else if (_T_53) begin
          lo <= rob_io_deq_bits_lo;
        end else if (_T_51) begin
          lo <= rob_io_deq_bits_lo;
        end else if (_T_49) begin
          lo <= rob_io_deq_bits_lo;
        end else if (_T_47) begin
          lo <= _T_30[31:0];
        end else if (_T_45) begin
          lo <= _T_30[31:0];
        end else if (_T_43) begin
          lo <= _T_36[31:0];
        end else if (_T_41) begin
          lo <= _T_36[31:0];
        end else begin
          lo <= 32'h0;
        end
      end
    end
    if (reset) begin
      mduid <= 6'h0;
    end else if (_T_7) begin
      mduid <= _T_9;
    end
  end
endmodule
module MSUPipelineStage(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input         io_fu_in_bits_wb_v,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_wen,
  input  [31:0] io_fu_in_bits_wb_data,
  input         io_fu_in_bits_wb_ip7,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  output        io_fu_out_valid,
  output        io_fu_out_bits_v,
  output [7:0]  io_fu_out_bits_id,
  output [31:0] io_fu_out_bits_pc,
  output [5:0]  io_fu_out_bits_instr_op,
  output [4:0]  io_fu_out_bits_instr_rs_idx,
  output [4:0]  io_fu_out_bits_instr_rt_idx,
  output [4:0]  io_fu_out_bits_instr_rd_idx,
  output [4:0]  io_fu_out_bits_instr_shamt,
  output [5:0]  io_fu_out_bits_instr_func,
  output [4:0]  io_fu_out_bits_rd_idx,
  output        io_fu_out_bits_wen,
  output [31:0] io_fu_out_bits_data,
  output        io_fu_out_bits_ip7,
  output        io_fu_out_bits_is_ds,
  output        io_fu_out_bits_is_br,
  output [31:0] io_fu_out_bits_npc
);
  wire  _T = io_fu_in_ready & io_fu_in_valid; // @[Decoupled.scala 40:37]
  reg  fu_in_wb_v; // @[Reg.scala 27:20]
  reg [31:0] _RAND_0;
  reg [7:0] fu_in_wb_id; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [31:0] fu_in_wb_pc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  reg [5:0] fu_in_wb_instr_op; // @[Reg.scala 27:20]
  reg [31:0] _RAND_3;
  reg [4:0] fu_in_wb_instr_rs_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [4:0] fu_in_wb_instr_rt_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [4:0] fu_in_wb_instr_rd_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [4:0] fu_in_wb_instr_shamt; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [5:0] fu_in_wb_instr_func; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  reg [4:0] fu_in_wb_rd_idx; // @[Reg.scala 27:20]
  reg [31:0] _RAND_9;
  reg  fu_in_wb_wen; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg [31:0] fu_in_wb_data; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg  fu_in_wb_ip7; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg  fu_in_wb_is_ds; // @[Reg.scala 27:20]
  reg [31:0] _RAND_13;
  reg  fu_in_wb_is_br; // @[Reg.scala 27:20]
  reg [31:0] _RAND_14;
  reg [31:0] fu_in_wb_npc; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  reg  fu_valid; // @[msu.scala 23:25]
  reg [31:0] _RAND_16;
  wire  _T_3 = ~_T; // @[msu.scala 27:9]
  wire  _T_4 = _T_3 & io_fu_out_valid; // @[msu.scala 27:26]
  wire  _GEN_17 = _T | fu_valid; // @[msu.scala 29:32]
  assign io_fu_in_ready = 1'h1; // @[msu.scala 24:18]
  assign io_fu_out_valid = fu_valid; // @[msu.scala 25:19]
  assign io_fu_out_bits_v = fu_in_wb_v; // @[msu.scala 26:18]
  assign io_fu_out_bits_id = fu_in_wb_id; // @[msu.scala 26:18]
  assign io_fu_out_bits_pc = fu_in_wb_pc; // @[msu.scala 26:18]
  assign io_fu_out_bits_instr_op = fu_in_wb_instr_op; // @[msu.scala 26:18]
  assign io_fu_out_bits_instr_rs_idx = fu_in_wb_instr_rs_idx; // @[msu.scala 26:18]
  assign io_fu_out_bits_instr_rt_idx = fu_in_wb_instr_rt_idx; // @[msu.scala 26:18]
  assign io_fu_out_bits_instr_rd_idx = fu_in_wb_instr_rd_idx; // @[msu.scala 26:18]
  assign io_fu_out_bits_instr_shamt = fu_in_wb_instr_shamt; // @[msu.scala 26:18]
  assign io_fu_out_bits_instr_func = fu_in_wb_instr_func; // @[msu.scala 26:18]
  assign io_fu_out_bits_rd_idx = fu_in_wb_rd_idx; // @[msu.scala 26:18]
  assign io_fu_out_bits_wen = fu_in_wb_wen; // @[msu.scala 26:18]
  assign io_fu_out_bits_data = fu_in_wb_data; // @[msu.scala 26:18]
  assign io_fu_out_bits_ip7 = fu_in_wb_ip7; // @[msu.scala 26:18]
  assign io_fu_out_bits_is_ds = fu_in_wb_is_ds; // @[msu.scala 26:18]
  assign io_fu_out_bits_is_br = fu_in_wb_is_br; // @[msu.scala 26:18]
  assign io_fu_out_bits_npc = fu_in_wb_npc; // @[msu.scala 26:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fu_in_wb_v = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  fu_in_wb_id = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  fu_in_wb_pc = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  fu_in_wb_instr_op = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  fu_in_wb_instr_rs_idx = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  fu_in_wb_instr_rt_idx = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fu_in_wb_instr_rd_idx = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  fu_in_wb_instr_shamt = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  fu_in_wb_instr_func = _RAND_8[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fu_in_wb_rd_idx = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fu_in_wb_wen = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fu_in_wb_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fu_in_wb_ip7 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fu_in_wb_is_ds = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fu_in_wb_is_br = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fu_in_wb_npc = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  fu_valid = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      fu_in_wb_v <= 1'h0;
    end else if (_T) begin
      fu_in_wb_v <= io_fu_in_bits_wb_v;
    end
    if (reset) begin
      fu_in_wb_id <= 8'h0;
    end else if (_T) begin
      fu_in_wb_id <= io_fu_in_bits_wb_id;
    end
    if (reset) begin
      fu_in_wb_pc <= 32'h0;
    end else if (_T) begin
      fu_in_wb_pc <= io_fu_in_bits_wb_pc;
    end
    if (reset) begin
      fu_in_wb_instr_op <= 6'h0;
    end else if (_T) begin
      fu_in_wb_instr_op <= io_fu_in_bits_wb_instr_op;
    end
    if (reset) begin
      fu_in_wb_instr_rs_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rs_idx <= io_fu_in_bits_wb_instr_rs_idx;
    end
    if (reset) begin
      fu_in_wb_instr_rt_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rt_idx <= io_fu_in_bits_wb_instr_rt_idx;
    end
    if (reset) begin
      fu_in_wb_instr_rd_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_rd_idx <= io_fu_in_bits_wb_instr_rd_idx;
    end
    if (reset) begin
      fu_in_wb_instr_shamt <= 5'h0;
    end else if (_T) begin
      fu_in_wb_instr_shamt <= io_fu_in_bits_wb_instr_shamt;
    end
    if (reset) begin
      fu_in_wb_instr_func <= 6'h0;
    end else if (_T) begin
      fu_in_wb_instr_func <= io_fu_in_bits_wb_instr_func;
    end
    if (reset) begin
      fu_in_wb_rd_idx <= 5'h0;
    end else if (_T) begin
      fu_in_wb_rd_idx <= io_fu_in_bits_wb_rd_idx;
    end
    if (reset) begin
      fu_in_wb_wen <= 1'h0;
    end else if (_T) begin
      fu_in_wb_wen <= io_fu_in_bits_wb_wen;
    end
    if (reset) begin
      fu_in_wb_data <= 32'h0;
    end else if (_T) begin
      fu_in_wb_data <= io_fu_in_bits_wb_data;
    end
    if (reset) begin
      fu_in_wb_ip7 <= 1'h0;
    end else if (_T) begin
      fu_in_wb_ip7 <= io_fu_in_bits_wb_ip7;
    end
    if (reset) begin
      fu_in_wb_is_ds <= 1'h0;
    end else if (_T) begin
      fu_in_wb_is_ds <= io_fu_in_bits_wb_is_ds;
    end
    if (reset) begin
      fu_in_wb_is_br <= 1'h0;
    end else if (_T) begin
      fu_in_wb_is_br <= io_fu_in_bits_wb_is_br;
    end
    if (reset) begin
      fu_in_wb_npc <= 32'h0;
    end else if (_T) begin
      fu_in_wb_npc <= io_fu_in_bits_wb_npc;
    end
    if (reset) begin
      fu_valid <= 1'h0;
    end else if (_T_4) begin
      fu_valid <= 1'h0;
    end else begin
      fu_valid <= _GEN_17;
    end
  end
endmodule
module MSU(
  input         clock,
  input         reset,
  output        io_fu_in_ready,
  input         io_fu_in_valid,
  input         io_fu_in_bits_wb_v,
  input  [7:0]  io_fu_in_bits_wb_id,
  input  [31:0] io_fu_in_bits_wb_pc,
  input  [5:0]  io_fu_in_bits_wb_instr_op,
  input  [4:0]  io_fu_in_bits_wb_instr_rs_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rt_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_rd_idx,
  input  [4:0]  io_fu_in_bits_wb_instr_shamt,
  input  [5:0]  io_fu_in_bits_wb_instr_func,
  input  [4:0]  io_fu_in_bits_wb_rd_idx,
  input         io_fu_in_bits_wb_wen,
  input  [31:0] io_fu_in_bits_wb_data,
  input         io_fu_in_bits_wb_ip7,
  input         io_fu_in_bits_wb_is_ds,
  input         io_fu_in_bits_wb_is_br,
  input  [31:0] io_fu_in_bits_wb_npc,
  input  [2:0]  io_fu_in_bits_ops_fu_type,
  input  [4:0]  io_fu_in_bits_ops_fu_op,
  input  [31:0] io_fu_in_bits_ops_op1,
  input  [31:0] io_fu_in_bits_ops_op2,
  input         io_fu_in_bits_is_cached,
  output        io_wb_valid,
  output        io_wb_bits_v,
  output [7:0]  io_wb_bits_id,
  output [31:0] io_wb_bits_pc,
  output [5:0]  io_wb_bits_instr_op,
  output [4:0]  io_wb_bits_instr_rs_idx,
  output [4:0]  io_wb_bits_instr_rt_idx,
  output [4:0]  io_wb_bits_instr_rd_idx,
  output [4:0]  io_wb_bits_instr_shamt,
  output [5:0]  io_wb_bits_instr_func,
  output [4:0]  io_wb_bits_rd_idx,
  output        io_wb_bits_wen,
  output [31:0] io_wb_bits_data,
  output        io_wb_bits_ip7,
  output        io_divider_data_dividend_tvalid,
  output        io_divider_data_divisor_tvalid,
  input         io_divider_data_dout_tvalid,
  output [39:0] io_divider_data_dividend_tdata,
  output [39:0] io_divider_data_divisor_tdata,
  input  [79:0] io_divider_data_dout_tdata,
  output [32:0] io_multiplier_data_a,
  output [32:0] io_multiplier_data_b,
  input  [65:0] io_multiplier_data_dout,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output        io_dmem_req_bits_is_cached,
  output [31:0] io_dmem_req_bits_addr,
  output [1:0]  io_dmem_req_bits_len,
  output [3:0]  io_dmem_req_bits_strb,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_func,
  input         io_dmem_resp_valid,
  input  [31:0] io_dmem_resp_bits_data
);
  wire  lsu_clock; // @[msu.scala 54:19]
  wire  lsu_reset; // @[msu.scala 54:19]
  wire  lsu_io_dmem_req_ready; // @[msu.scala 54:19]
  wire  lsu_io_dmem_req_valid; // @[msu.scala 54:19]
  wire  lsu_io_dmem_req_bits_is_cached; // @[msu.scala 54:19]
  wire [31:0] lsu_io_dmem_req_bits_addr; // @[msu.scala 54:19]
  wire [1:0] lsu_io_dmem_req_bits_len; // @[msu.scala 54:19]
  wire [3:0] lsu_io_dmem_req_bits_strb; // @[msu.scala 54:19]
  wire [31:0] lsu_io_dmem_req_bits_data; // @[msu.scala 54:19]
  wire  lsu_io_dmem_req_bits_func; // @[msu.scala 54:19]
  wire  lsu_io_dmem_resp_ready; // @[msu.scala 54:19]
  wire  lsu_io_dmem_resp_valid; // @[msu.scala 54:19]
  wire [31:0] lsu_io_dmem_resp_bits_data; // @[msu.scala 54:19]
  wire  lsu_io_fu_in_ready; // @[msu.scala 54:19]
  wire  lsu_io_fu_in_valid; // @[msu.scala 54:19]
  wire [7:0] lsu_io_fu_in_bits_wb_id; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_in_bits_wb_pc; // @[msu.scala 54:19]
  wire [5:0] lsu_io_fu_in_bits_wb_instr_op; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_in_bits_wb_instr_rs_idx; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_in_bits_wb_instr_rt_idx; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_in_bits_wb_instr_rd_idx; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_in_bits_wb_instr_shamt; // @[msu.scala 54:19]
  wire [5:0] lsu_io_fu_in_bits_wb_instr_func; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_in_bits_wb_rd_idx; // @[msu.scala 54:19]
  wire  lsu_io_fu_in_bits_wb_ip7; // @[msu.scala 54:19]
  wire  lsu_io_fu_in_bits_wb_is_br; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_in_bits_wb_npc; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_in_bits_ops_fu_op; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_in_bits_ops_op1; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_in_bits_ops_op2; // @[msu.scala 54:19]
  wire  lsu_io_fu_in_bits_is_cached; // @[msu.scala 54:19]
  wire  lsu_io_fu_out_valid; // @[msu.scala 54:19]
  wire  lsu_io_fu_out_bits_v; // @[msu.scala 54:19]
  wire [7:0] lsu_io_fu_out_bits_id; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_out_bits_pc; // @[msu.scala 54:19]
  wire [5:0] lsu_io_fu_out_bits_instr_op; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_out_bits_instr_rs_idx; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_out_bits_instr_rt_idx; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_out_bits_instr_rd_idx; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_out_bits_instr_shamt; // @[msu.scala 54:19]
  wire [5:0] lsu_io_fu_out_bits_instr_func; // @[msu.scala 54:19]
  wire [4:0] lsu_io_fu_out_bits_rd_idx; // @[msu.scala 54:19]
  wire  lsu_io_fu_out_bits_wen; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_out_bits_data; // @[msu.scala 54:19]
  wire  lsu_io_fu_out_bits_ip7; // @[msu.scala 54:19]
  wire  lsu_io_fu_out_bits_is_br; // @[msu.scala 54:19]
  wire [31:0] lsu_io_fu_out_bits_npc; // @[msu.scala 54:19]
  wire  lsu_io_working; // @[msu.scala 54:19]
  wire  mdu_clock; // @[msu.scala 55:19]
  wire  mdu_reset; // @[msu.scala 55:19]
  wire  mdu_io_fu_in_ready; // @[msu.scala 55:19]
  wire  mdu_io_fu_in_valid; // @[msu.scala 55:19]
  wire [7:0] mdu_io_fu_in_bits_wb_id; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_in_bits_wb_pc; // @[msu.scala 55:19]
  wire [5:0] mdu_io_fu_in_bits_wb_instr_op; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_in_bits_wb_instr_rs_idx; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_in_bits_wb_instr_rt_idx; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_in_bits_wb_instr_rd_idx; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_in_bits_wb_instr_shamt; // @[msu.scala 55:19]
  wire [5:0] mdu_io_fu_in_bits_wb_instr_func; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_in_bits_wb_rd_idx; // @[msu.scala 55:19]
  wire  mdu_io_fu_in_bits_wb_ip7; // @[msu.scala 55:19]
  wire  mdu_io_fu_in_bits_wb_is_ds; // @[msu.scala 55:19]
  wire  mdu_io_fu_in_bits_wb_is_br; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_in_bits_wb_npc; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_in_bits_ops_fu_op; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_in_bits_ops_op1; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_in_bits_ops_op2; // @[msu.scala 55:19]
  wire  mdu_io_fu_out_valid; // @[msu.scala 55:19]
  wire  mdu_io_fu_out_bits_v; // @[msu.scala 55:19]
  wire [7:0] mdu_io_fu_out_bits_id; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_out_bits_pc; // @[msu.scala 55:19]
  wire [5:0] mdu_io_fu_out_bits_instr_op; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_out_bits_instr_rs_idx; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_out_bits_instr_rt_idx; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_out_bits_instr_rd_idx; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_out_bits_instr_shamt; // @[msu.scala 55:19]
  wire [5:0] mdu_io_fu_out_bits_instr_func; // @[msu.scala 55:19]
  wire [4:0] mdu_io_fu_out_bits_rd_idx; // @[msu.scala 55:19]
  wire  mdu_io_fu_out_bits_wen; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_out_bits_data; // @[msu.scala 55:19]
  wire  mdu_io_fu_out_bits_ip7; // @[msu.scala 55:19]
  wire  mdu_io_fu_out_bits_is_ds; // @[msu.scala 55:19]
  wire  mdu_io_fu_out_bits_is_br; // @[msu.scala 55:19]
  wire [31:0] mdu_io_fu_out_bits_npc; // @[msu.scala 55:19]
  wire  mdu_io_working; // @[msu.scala 55:19]
  wire  mdu_io_divider_data_dividend_tvalid; // @[msu.scala 55:19]
  wire  mdu_io_divider_data_divisor_tvalid; // @[msu.scala 55:19]
  wire  mdu_io_divider_data_dout_tvalid; // @[msu.scala 55:19]
  wire [39:0] mdu_io_divider_data_dividend_tdata; // @[msu.scala 55:19]
  wire [39:0] mdu_io_divider_data_divisor_tdata; // @[msu.scala 55:19]
  wire [79:0] mdu_io_divider_data_dout_tdata; // @[msu.scala 55:19]
  wire [32:0] mdu_io_multiplier_data_a; // @[msu.scala 55:19]
  wire [32:0] mdu_io_multiplier_data_b; // @[msu.scala 55:19]
  wire [65:0] mdu_io_multiplier_data_dout; // @[msu.scala 55:19]
  wire  psu_clock; // @[msu.scala 56:19]
  wire  psu_reset; // @[msu.scala 56:19]
  wire  psu_io_fu_in_ready; // @[msu.scala 56:19]
  wire  psu_io_fu_in_valid; // @[msu.scala 56:19]
  wire  psu_io_fu_in_bits_wb_v; // @[msu.scala 56:19]
  wire [7:0] psu_io_fu_in_bits_wb_id; // @[msu.scala 56:19]
  wire [31:0] psu_io_fu_in_bits_wb_pc; // @[msu.scala 56:19]
  wire [5:0] psu_io_fu_in_bits_wb_instr_op; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_in_bits_wb_instr_rs_idx; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_in_bits_wb_instr_rt_idx; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_in_bits_wb_instr_rd_idx; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_in_bits_wb_instr_shamt; // @[msu.scala 56:19]
  wire [5:0] psu_io_fu_in_bits_wb_instr_func; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_in_bits_wb_rd_idx; // @[msu.scala 56:19]
  wire  psu_io_fu_in_bits_wb_wen; // @[msu.scala 56:19]
  wire [31:0] psu_io_fu_in_bits_wb_data; // @[msu.scala 56:19]
  wire  psu_io_fu_in_bits_wb_ip7; // @[msu.scala 56:19]
  wire  psu_io_fu_in_bits_wb_is_ds; // @[msu.scala 56:19]
  wire  psu_io_fu_in_bits_wb_is_br; // @[msu.scala 56:19]
  wire [31:0] psu_io_fu_in_bits_wb_npc; // @[msu.scala 56:19]
  wire  psu_io_fu_out_valid; // @[msu.scala 56:19]
  wire  psu_io_fu_out_bits_v; // @[msu.scala 56:19]
  wire [7:0] psu_io_fu_out_bits_id; // @[msu.scala 56:19]
  wire [31:0] psu_io_fu_out_bits_pc; // @[msu.scala 56:19]
  wire [5:0] psu_io_fu_out_bits_instr_op; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_out_bits_instr_rs_idx; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_out_bits_instr_rt_idx; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_out_bits_instr_rd_idx; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_out_bits_instr_shamt; // @[msu.scala 56:19]
  wire [5:0] psu_io_fu_out_bits_instr_func; // @[msu.scala 56:19]
  wire [4:0] psu_io_fu_out_bits_rd_idx; // @[msu.scala 56:19]
  wire  psu_io_fu_out_bits_wen; // @[msu.scala 56:19]
  wire [31:0] psu_io_fu_out_bits_data; // @[msu.scala 56:19]
  wire  psu_io_fu_out_bits_ip7; // @[msu.scala 56:19]
  wire  psu_io_fu_out_bits_is_ds; // @[msu.scala 56:19]
  wire  psu_io_fu_out_bits_is_br; // @[msu.scala 56:19]
  wire [31:0] psu_io_fu_out_bits_npc; // @[msu.scala 56:19]
  wire  _T = ~mdu_io_working; // @[msu.scala 59:16]
  wire  _T_1 = io_fu_in_bits_ops_fu_type == 3'h3; // @[msu.scala 60:31]
  wire  to_lsu = _T & _T_1; // @[msu.scala 59:32]
  wire  _T_3 = ~lsu_io_working; // @[msu.scala 67:16]
  wire  _T_4 = io_fu_in_bits_ops_fu_type == 3'h4; // @[msu.scala 68:31]
  wire  to_mdu = _T_3 & _T_4; // @[msu.scala 67:32]
  wire  _T_8 = _T_3 & _T; // @[msu.scala 76:32]
  wire  _T_9 = io_fu_in_bits_ops_fu_type != 3'h3; // @[msu.scala 77:32]
  wire  _T_10 = io_fu_in_bits_ops_fu_type != 3'h4; // @[msu.scala 78:31]
  wire  _T_11 = _T_9 & _T_10; // @[msu.scala 77:43]
  wire  to_psu = _T_8 & _T_11; // @[msu.scala 76:51]
  wire  _T_19 = ~io_fu_in_bits_ops_fu_op[3]; // @[msu.scala 80:54]
  wire  is_lsu_load = _T_1 & _T_19; // @[msu.scala 79:58]
  wire  _T_22 = to_lsu & lsu_io_fu_in_ready; // @[msu.scala 88:29]
  wire  _T_24 = _T_22 | to_mdu; // @[msu.scala 88:52]
  wire  _T_27 = lsu_io_fu_out_valid | mdu_io_fu_out_valid; // @[msu.scala 91:38]
  wire [78:0] _T_35 = {lsu_io_fu_out_bits_instr_func,lsu_io_fu_out_bits_rd_idx,lsu_io_fu_out_bits_wen,lsu_io_fu_out_bits_data,lsu_io_fu_out_bits_ip7,1'h0,lsu_io_fu_out_bits_is_br,lsu_io_fu_out_bits_npc}; // @[Mux.scala 27:72]
  wire [145:0] _T_43 = {lsu_io_fu_out_bits_v,lsu_io_fu_out_bits_id,lsu_io_fu_out_bits_pc,lsu_io_fu_out_bits_instr_op,lsu_io_fu_out_bits_instr_rs_idx,lsu_io_fu_out_bits_instr_rt_idx,lsu_io_fu_out_bits_instr_rd_idx,lsu_io_fu_out_bits_instr_shamt,_T_35}; // @[Mux.scala 27:72]
  wire [145:0] _T_44 = lsu_io_fu_out_valid ? _T_43 : 146'h0; // @[Mux.scala 27:72]
  wire [78:0] _T_51 = {mdu_io_fu_out_bits_instr_func,mdu_io_fu_out_bits_rd_idx,mdu_io_fu_out_bits_wen,mdu_io_fu_out_bits_data,mdu_io_fu_out_bits_ip7,mdu_io_fu_out_bits_is_ds,mdu_io_fu_out_bits_is_br,mdu_io_fu_out_bits_npc}; // @[Mux.scala 27:72]
  wire [145:0] _T_59 = {mdu_io_fu_out_bits_v,mdu_io_fu_out_bits_id,mdu_io_fu_out_bits_pc,mdu_io_fu_out_bits_instr_op,mdu_io_fu_out_bits_instr_rs_idx,mdu_io_fu_out_bits_instr_rt_idx,mdu_io_fu_out_bits_instr_rd_idx,mdu_io_fu_out_bits_instr_shamt,_T_51}; // @[Mux.scala 27:72]
  wire [145:0] _T_60 = mdu_io_fu_out_valid ? _T_59 : 146'h0; // @[Mux.scala 27:72]
  wire [78:0] _T_67 = {psu_io_fu_out_bits_instr_func,psu_io_fu_out_bits_rd_idx,psu_io_fu_out_bits_wen,psu_io_fu_out_bits_data,psu_io_fu_out_bits_ip7,psu_io_fu_out_bits_is_ds,psu_io_fu_out_bits_is_br,psu_io_fu_out_bits_npc}; // @[Mux.scala 27:72]
  wire [145:0] _T_75 = {psu_io_fu_out_bits_v,psu_io_fu_out_bits_id,psu_io_fu_out_bits_pc,psu_io_fu_out_bits_instr_op,psu_io_fu_out_bits_instr_rs_idx,psu_io_fu_out_bits_instr_rt_idx,psu_io_fu_out_bits_instr_rd_idx,psu_io_fu_out_bits_instr_shamt,_T_67}; // @[Mux.scala 27:72]
  wire [145:0] _T_76 = psu_io_fu_out_valid ? _T_75 : 146'h0; // @[Mux.scala 27:72]
  wire [145:0] _T_77 = _T_44 | _T_60; // @[Mux.scala 27:72]
  wire [145:0] _T_78 = _T_77 | _T_76; // @[Mux.scala 27:72]
  wire [2:0] _T_98 = {lsu_io_fu_out_valid,mdu_io_fu_out_valid,psu_io_fu_out_valid}; // @[Cat.scala 29:58]
  wire  _T_99 = _T_98 != 3'h0; // @[utils.scala 129:38]
  wire  _T_100 = ~_T_99; // @[utils.scala 129:27]
  wire  _T_101 = lsu_io_fu_out_valid; // @[utils.scala 123:35]
  wire  _T_102 = ~mdu_io_fu_out_valid; // @[utils.scala 123:44]
  wire  _T_103 = ~psu_io_fu_out_valid; // @[utils.scala 123:44]
  wire [2:0] _T_105 = {_T_101,_T_102,_T_103}; // @[Cat.scala 29:58]
  wire  _T_106 = _T_105 == 3'h7; // @[utils.scala 123:63]
  wire  _T_107 = ~lsu_io_fu_out_valid; // @[utils.scala 123:44]
  wire  _T_108 = mdu_io_fu_out_valid; // @[utils.scala 123:35]
  wire [2:0] _T_111 = {_T_107,_T_108,_T_103}; // @[Cat.scala 29:58]
  wire  _T_112 = _T_111 == 3'h7; // @[utils.scala 123:63]
  wire  _T_115 = psu_io_fu_out_valid; // @[utils.scala 123:35]
  wire [2:0] _T_117 = {_T_107,_T_102,_T_115}; // @[Cat.scala 29:58]
  wire  _T_118 = _T_117 == 3'h7; // @[utils.scala 123:63]
  wire [2:0] _T_120 = {_T_106,_T_112,_T_118}; // @[Cat.scala 29:58]
  wire  _T_121 = _T_120 != 3'h0; // @[utils.scala 124:9]
  reg  _T_123; // @[msu.scala 108:18]
  reg [31:0] _RAND_0;
  reg [30:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_1;
  wire  _T_125 = value == 31'h7ffffffe; // @[Counter.scala 38:24]
  wire [30:0] _T_127 = value + 31'h1; // @[Counter.scala 39:22]
  wire  _T_129 = _T_123 | reset; // @[msu.scala 108:10]
  wire  _T_130 = ~_T_129; // @[msu.scala 108:10]
  LSU lsu ( // @[msu.scala 54:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_dmem_req_ready(lsu_io_dmem_req_ready),
    .io_dmem_req_valid(lsu_io_dmem_req_valid),
    .io_dmem_req_bits_is_cached(lsu_io_dmem_req_bits_is_cached),
    .io_dmem_req_bits_addr(lsu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_len(lsu_io_dmem_req_bits_len),
    .io_dmem_req_bits_strb(lsu_io_dmem_req_bits_strb),
    .io_dmem_req_bits_data(lsu_io_dmem_req_bits_data),
    .io_dmem_req_bits_func(lsu_io_dmem_req_bits_func),
    .io_dmem_resp_ready(lsu_io_dmem_resp_ready),
    .io_dmem_resp_valid(lsu_io_dmem_resp_valid),
    .io_dmem_resp_bits_data(lsu_io_dmem_resp_bits_data),
    .io_fu_in_ready(lsu_io_fu_in_ready),
    .io_fu_in_valid(lsu_io_fu_in_valid),
    .io_fu_in_bits_wb_id(lsu_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(lsu_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(lsu_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(lsu_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(lsu_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(lsu_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(lsu_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(lsu_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(lsu_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_ip7(lsu_io_fu_in_bits_wb_ip7),
    .io_fu_in_bits_wb_is_br(lsu_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(lsu_io_fu_in_bits_wb_npc),
    .io_fu_in_bits_ops_fu_op(lsu_io_fu_in_bits_ops_fu_op),
    .io_fu_in_bits_ops_op1(lsu_io_fu_in_bits_ops_op1),
    .io_fu_in_bits_ops_op2(lsu_io_fu_in_bits_ops_op2),
    .io_fu_in_bits_is_cached(lsu_io_fu_in_bits_is_cached),
    .io_fu_out_valid(lsu_io_fu_out_valid),
    .io_fu_out_bits_v(lsu_io_fu_out_bits_v),
    .io_fu_out_bits_id(lsu_io_fu_out_bits_id),
    .io_fu_out_bits_pc(lsu_io_fu_out_bits_pc),
    .io_fu_out_bits_instr_op(lsu_io_fu_out_bits_instr_op),
    .io_fu_out_bits_instr_rs_idx(lsu_io_fu_out_bits_instr_rs_idx),
    .io_fu_out_bits_instr_rt_idx(lsu_io_fu_out_bits_instr_rt_idx),
    .io_fu_out_bits_instr_rd_idx(lsu_io_fu_out_bits_instr_rd_idx),
    .io_fu_out_bits_instr_shamt(lsu_io_fu_out_bits_instr_shamt),
    .io_fu_out_bits_instr_func(lsu_io_fu_out_bits_instr_func),
    .io_fu_out_bits_rd_idx(lsu_io_fu_out_bits_rd_idx),
    .io_fu_out_bits_wen(lsu_io_fu_out_bits_wen),
    .io_fu_out_bits_data(lsu_io_fu_out_bits_data),
    .io_fu_out_bits_ip7(lsu_io_fu_out_bits_ip7),
    .io_fu_out_bits_is_br(lsu_io_fu_out_bits_is_br),
    .io_fu_out_bits_npc(lsu_io_fu_out_bits_npc),
    .io_working(lsu_io_working)
  );
  MDU mdu ( // @[msu.scala 55:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_fu_in_ready(mdu_io_fu_in_ready),
    .io_fu_in_valid(mdu_io_fu_in_valid),
    .io_fu_in_bits_wb_id(mdu_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(mdu_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(mdu_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(mdu_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(mdu_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(mdu_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(mdu_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(mdu_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(mdu_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_ip7(mdu_io_fu_in_bits_wb_ip7),
    .io_fu_in_bits_wb_is_ds(mdu_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(mdu_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(mdu_io_fu_in_bits_wb_npc),
    .io_fu_in_bits_ops_fu_op(mdu_io_fu_in_bits_ops_fu_op),
    .io_fu_in_bits_ops_op1(mdu_io_fu_in_bits_ops_op1),
    .io_fu_in_bits_ops_op2(mdu_io_fu_in_bits_ops_op2),
    .io_fu_out_valid(mdu_io_fu_out_valid),
    .io_fu_out_bits_v(mdu_io_fu_out_bits_v),
    .io_fu_out_bits_id(mdu_io_fu_out_bits_id),
    .io_fu_out_bits_pc(mdu_io_fu_out_bits_pc),
    .io_fu_out_bits_instr_op(mdu_io_fu_out_bits_instr_op),
    .io_fu_out_bits_instr_rs_idx(mdu_io_fu_out_bits_instr_rs_idx),
    .io_fu_out_bits_instr_rt_idx(mdu_io_fu_out_bits_instr_rt_idx),
    .io_fu_out_bits_instr_rd_idx(mdu_io_fu_out_bits_instr_rd_idx),
    .io_fu_out_bits_instr_shamt(mdu_io_fu_out_bits_instr_shamt),
    .io_fu_out_bits_instr_func(mdu_io_fu_out_bits_instr_func),
    .io_fu_out_bits_rd_idx(mdu_io_fu_out_bits_rd_idx),
    .io_fu_out_bits_wen(mdu_io_fu_out_bits_wen),
    .io_fu_out_bits_data(mdu_io_fu_out_bits_data),
    .io_fu_out_bits_ip7(mdu_io_fu_out_bits_ip7),
    .io_fu_out_bits_is_ds(mdu_io_fu_out_bits_is_ds),
    .io_fu_out_bits_is_br(mdu_io_fu_out_bits_is_br),
    .io_fu_out_bits_npc(mdu_io_fu_out_bits_npc),
    .io_working(mdu_io_working),
    .io_divider_data_dividend_tvalid(mdu_io_divider_data_dividend_tvalid),
    .io_divider_data_divisor_tvalid(mdu_io_divider_data_divisor_tvalid),
    .io_divider_data_dout_tvalid(mdu_io_divider_data_dout_tvalid),
    .io_divider_data_dividend_tdata(mdu_io_divider_data_dividend_tdata),
    .io_divider_data_divisor_tdata(mdu_io_divider_data_divisor_tdata),
    .io_divider_data_dout_tdata(mdu_io_divider_data_dout_tdata),
    .io_multiplier_data_a(mdu_io_multiplier_data_a),
    .io_multiplier_data_b(mdu_io_multiplier_data_b),
    .io_multiplier_data_dout(mdu_io_multiplier_data_dout)
  );
  MSUPipelineStage psu ( // @[msu.scala 56:19]
    .clock(psu_clock),
    .reset(psu_reset),
    .io_fu_in_ready(psu_io_fu_in_ready),
    .io_fu_in_valid(psu_io_fu_in_valid),
    .io_fu_in_bits_wb_v(psu_io_fu_in_bits_wb_v),
    .io_fu_in_bits_wb_id(psu_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(psu_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(psu_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(psu_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(psu_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(psu_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(psu_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(psu_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(psu_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_wen(psu_io_fu_in_bits_wb_wen),
    .io_fu_in_bits_wb_data(psu_io_fu_in_bits_wb_data),
    .io_fu_in_bits_wb_ip7(psu_io_fu_in_bits_wb_ip7),
    .io_fu_in_bits_wb_is_ds(psu_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(psu_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(psu_io_fu_in_bits_wb_npc),
    .io_fu_out_valid(psu_io_fu_out_valid),
    .io_fu_out_bits_v(psu_io_fu_out_bits_v),
    .io_fu_out_bits_id(psu_io_fu_out_bits_id),
    .io_fu_out_bits_pc(psu_io_fu_out_bits_pc),
    .io_fu_out_bits_instr_op(psu_io_fu_out_bits_instr_op),
    .io_fu_out_bits_instr_rs_idx(psu_io_fu_out_bits_instr_rs_idx),
    .io_fu_out_bits_instr_rt_idx(psu_io_fu_out_bits_instr_rt_idx),
    .io_fu_out_bits_instr_rd_idx(psu_io_fu_out_bits_instr_rd_idx),
    .io_fu_out_bits_instr_shamt(psu_io_fu_out_bits_instr_shamt),
    .io_fu_out_bits_instr_func(psu_io_fu_out_bits_instr_func),
    .io_fu_out_bits_rd_idx(psu_io_fu_out_bits_rd_idx),
    .io_fu_out_bits_wen(psu_io_fu_out_bits_wen),
    .io_fu_out_bits_data(psu_io_fu_out_bits_data),
    .io_fu_out_bits_ip7(psu_io_fu_out_bits_ip7),
    .io_fu_out_bits_is_ds(psu_io_fu_out_bits_is_ds),
    .io_fu_out_bits_is_br(psu_io_fu_out_bits_is_br),
    .io_fu_out_bits_npc(psu_io_fu_out_bits_npc)
  );
  assign io_fu_in_ready = _T_24 | to_psu; // @[msu.scala 88:18]
  assign io_wb_valid = _T_27 | psu_io_fu_out_valid; // @[msu.scala 91:15]
  assign io_wb_bits_v = _T_78[145]; // @[msu.scala 92:14]
  assign io_wb_bits_id = _T_78[144:137]; // @[msu.scala 92:14]
  assign io_wb_bits_pc = _T_78[136:105]; // @[msu.scala 92:14]
  assign io_wb_bits_instr_op = _T_78[104:99]; // @[msu.scala 92:14]
  assign io_wb_bits_instr_rs_idx = _T_78[98:94]; // @[msu.scala 92:14]
  assign io_wb_bits_instr_rt_idx = _T_78[93:89]; // @[msu.scala 92:14]
  assign io_wb_bits_instr_rd_idx = _T_78[88:84]; // @[msu.scala 92:14]
  assign io_wb_bits_instr_shamt = _T_78[83:79]; // @[msu.scala 92:14]
  assign io_wb_bits_instr_func = _T_78[78:73]; // @[msu.scala 92:14]
  assign io_wb_bits_rd_idx = _T_78[72:68]; // @[msu.scala 92:14]
  assign io_wb_bits_wen = _T_78[67]; // @[msu.scala 92:14]
  assign io_wb_bits_data = _T_78[66:35]; // @[msu.scala 92:14]
  assign io_wb_bits_ip7 = _T_78[34]; // @[msu.scala 92:14]
  assign io_divider_data_dividend_tvalid = mdu_io_divider_data_dividend_tvalid; // @[msu.scala 71:18]
  assign io_divider_data_divisor_tvalid = mdu_io_divider_data_divisor_tvalid; // @[msu.scala 71:18]
  assign io_divider_data_dividend_tdata = mdu_io_divider_data_dividend_tdata; // @[msu.scala 71:18]
  assign io_divider_data_divisor_tdata = mdu_io_divider_data_divisor_tdata; // @[msu.scala 71:18]
  assign io_multiplier_data_a = mdu_io_multiplier_data_a; // @[msu.scala 72:21]
  assign io_multiplier_data_b = mdu_io_multiplier_data_b; // @[msu.scala 72:21]
  assign io_dmem_req_valid = lsu_io_dmem_req_valid; // @[msu.scala 63:15]
  assign io_dmem_req_bits_is_cached = lsu_io_dmem_req_bits_is_cached; // @[msu.scala 63:15]
  assign io_dmem_req_bits_addr = lsu_io_dmem_req_bits_addr; // @[msu.scala 63:15]
  assign io_dmem_req_bits_len = lsu_io_dmem_req_bits_len; // @[msu.scala 63:15]
  assign io_dmem_req_bits_strb = lsu_io_dmem_req_bits_strb; // @[msu.scala 63:15]
  assign io_dmem_req_bits_data = lsu_io_dmem_req_bits_data; // @[msu.scala 63:15]
  assign io_dmem_req_bits_func = lsu_io_dmem_req_bits_func; // @[msu.scala 63:15]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_dmem_req_ready = io_dmem_req_ready; // @[msu.scala 63:15]
  assign lsu_io_dmem_resp_valid = io_dmem_resp_valid; // @[msu.scala 63:15]
  assign lsu_io_dmem_resp_bits_data = io_dmem_resp_bits_data; // @[msu.scala 63:15]
  assign lsu_io_fu_in_valid = io_fu_in_valid & to_lsu; // @[msu.scala 61:22]
  assign lsu_io_fu_in_bits_wb_id = io_fu_in_bits_wb_id; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_pc = io_fu_in_bits_wb_pc; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_wb_npc = io_fu_in_bits_wb_npc; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_ops_fu_op = io_fu_in_bits_ops_fu_op; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_ops_op1 = io_fu_in_bits_ops_op1; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_ops_op2 = io_fu_in_bits_ops_op2; // @[msu.scala 62:21]
  assign lsu_io_fu_in_bits_is_cached = io_fu_in_bits_is_cached; // @[msu.scala 62:21]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_fu_in_valid = io_fu_in_valid & to_mdu; // @[msu.scala 69:22]
  assign mdu_io_fu_in_bits_wb_id = io_fu_in_bits_wb_id; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_pc = io_fu_in_bits_wb_pc; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_is_ds = io_fu_in_bits_wb_is_ds; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_wb_npc = io_fu_in_bits_wb_npc; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_ops_fu_op = io_fu_in_bits_ops_fu_op; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_ops_op1 = io_fu_in_bits_ops_op1; // @[msu.scala 70:21]
  assign mdu_io_fu_in_bits_ops_op2 = io_fu_in_bits_ops_op2; // @[msu.scala 70:21]
  assign mdu_io_divider_data_dout_tvalid = io_divider_data_dout_tvalid; // @[msu.scala 71:18]
  assign mdu_io_divider_data_dout_tdata = io_divider_data_dout_tdata; // @[msu.scala 71:18]
  assign mdu_io_multiplier_data_dout = io_multiplier_data_dout; // @[msu.scala 72:21]
  assign psu_clock = clock;
  assign psu_reset = reset;
  assign psu_io_fu_in_valid = io_fu_in_valid & to_psu; // @[msu.scala 81:22]
  assign psu_io_fu_in_bits_wb_v = is_lsu_load | io_fu_in_bits_wb_v; // @[msu.scala 82:24 msu.scala 83:26]
  assign psu_io_fu_in_bits_wb_id = io_fu_in_bits_wb_id; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_pc = io_fu_in_bits_wb_pc; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_instr_op = io_fu_in_bits_wb_instr_op; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_instr_rs_idx = io_fu_in_bits_wb_instr_rs_idx; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_instr_rt_idx = io_fu_in_bits_wb_instr_rt_idx; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_instr_rd_idx = io_fu_in_bits_wb_instr_rd_idx; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_instr_shamt = io_fu_in_bits_wb_instr_shamt; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_instr_func = io_fu_in_bits_wb_instr_func; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_rd_idx = io_fu_in_bits_wb_rd_idx; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_wen = io_fu_in_bits_wb_wen; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_data = io_fu_in_bits_wb_data; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_ip7 = io_fu_in_bits_wb_ip7; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_is_ds = io_fu_in_bits_wb_is_ds; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_is_br = io_fu_in_bits_wb_is_br; // @[msu.scala 82:24]
  assign psu_io_fu_in_bits_wb_npc = io_fu_in_bits_wb_npc; // @[msu.scala 82:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_123 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  value = _RAND_1[30:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_123 <= _T_100 | _T_121;
    if (reset) begin
      value <= 31'h0;
    end else if (_T_125) begin
      value <= 31'h0;
    end else begin
      value <= _T_127;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_130) begin
          $fwrite(32'h80000002,"Assertion failed: cycles: %d\n    at msu.scala:108 assert (RegNext(AtMost1H(lsu.io.fu_out.valid,\n",value); // @[msu.scala 108:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_130) begin
          $fatal; // @[msu.scala 108:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output        io_imem_req_bits_is_cached,
  output [31:0] io_imem_req_bits_addr,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [31:0] io_imem_resp_bits_data,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output        io_dmem_req_bits_is_cached,
  output [31:0] io_dmem_req_bits_addr,
  output [1:0]  io_dmem_req_bits_len,
  output [3:0]  io_dmem_req_bits_strb,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_func,
  input         io_dmem_resp_valid,
  input  [31:0] io_dmem_resp_bits_data,
  output        io_icache_control_valid,
  output [2:0]  io_icache_control_bits_op,
  output [31:0] io_icache_control_bits_addr,
  output        io_commit_valid,
  output [31:0] io_commit_pc,
  output [31:0] io_commit_instr,
  output        io_commit_ip7,
  output [31:0] io_commit_gpr_0,
  output [31:0] io_commit_gpr_1,
  output [31:0] io_commit_gpr_2,
  output [31:0] io_commit_gpr_3,
  output [31:0] io_commit_gpr_4,
  output [31:0] io_commit_gpr_5,
  output [31:0] io_commit_gpr_6,
  output [31:0] io_commit_gpr_7,
  output [31:0] io_commit_gpr_8,
  output [31:0] io_commit_gpr_9,
  output [31:0] io_commit_gpr_10,
  output [31:0] io_commit_gpr_11,
  output [31:0] io_commit_gpr_12,
  output [31:0] io_commit_gpr_13,
  output [31:0] io_commit_gpr_14,
  output [31:0] io_commit_gpr_15,
  output [31:0] io_commit_gpr_16,
  output [31:0] io_commit_gpr_17,
  output [31:0] io_commit_gpr_18,
  output [31:0] io_commit_gpr_19,
  output [31:0] io_commit_gpr_20,
  output [31:0] io_commit_gpr_21,
  output [31:0] io_commit_gpr_22,
  output [31:0] io_commit_gpr_23,
  output [31:0] io_commit_gpr_24,
  output [31:0] io_commit_gpr_25,
  output [31:0] io_commit_gpr_26,
  output [31:0] io_commit_gpr_27,
  output [31:0] io_commit_gpr_28,
  output [31:0] io_commit_gpr_29,
  output [31:0] io_commit_gpr_30,
  output [31:0] io_commit_gpr_31,
  output [4:0]  io_commit_rd_idx,
  output [31:0] io_commit_wdata,
  output        io_commit_wen,
  output        io_br_flush,
  output        io_ex_flush,
  output [32:0] io_multiplier_data_a,
  output [32:0] io_multiplier_data_b,
  input  [65:0] io_multiplier_data_dout,
  output        io_divider_data_dividend_tvalid,
  output        io_divider_data_divisor_tvalid,
  input         io_divider_data_dout_tvalid,
  output [39:0] io_divider_data_dividend_tdata,
  output [39:0] io_divider_data_divisor_tdata,
  input  [79:0] io_divider_data_dout_tdata
);
  wire  rf_clock; // @[core.scala 24:19]
  wire  rf_reset; // @[core.scala 24:19]
  wire  rf_io_bp_valid; // @[core.scala 24:19]
  wire  rf_io_bp_bits_v; // @[core.scala 24:19]
  wire [4:0] rf_io_bp_bits_rd_idx; // @[core.scala 24:19]
  wire  rf_io_bp_bits_wen; // @[core.scala 24:19]
  wire [31:0] rf_io_bp_bits_data; // @[core.scala 24:19]
  wire  rf_io_wb_valid; // @[core.scala 24:19]
  wire  rf_io_wb_bits_v; // @[core.scala 24:19]
  wire [7:0] rf_io_wb_bits_id; // @[core.scala 24:19]
  wire [31:0] rf_io_wb_bits_pc; // @[core.scala 24:19]
  wire [5:0] rf_io_wb_bits_instr_op; // @[core.scala 24:19]
  wire [4:0] rf_io_wb_bits_instr_rs_idx; // @[core.scala 24:19]
  wire [4:0] rf_io_wb_bits_instr_rt_idx; // @[core.scala 24:19]
  wire [4:0] rf_io_wb_bits_instr_rd_idx; // @[core.scala 24:19]
  wire [4:0] rf_io_wb_bits_instr_shamt; // @[core.scala 24:19]
  wire [5:0] rf_io_wb_bits_instr_func; // @[core.scala 24:19]
  wire [4:0] rf_io_wb_bits_rd_idx; // @[core.scala 24:19]
  wire  rf_io_wb_bits_wen; // @[core.scala 24:19]
  wire [31:0] rf_io_wb_bits_data; // @[core.scala 24:19]
  wire  rf_io_wb_bits_ip7; // @[core.scala 24:19]
  wire [4:0] rf_io_rfio_rs_idx; // @[core.scala 24:19]
  wire [4:0] rf_io_rfio_rt_idx; // @[core.scala 24:19]
  wire  rf_io_rfio_wen; // @[core.scala 24:19]
  wire [7:0] rf_io_rfio_wid; // @[core.scala 24:19]
  wire [4:0] rf_io_rfio_rd_idx; // @[core.scala 24:19]
  wire  rf_io_rfio_rs_data_valid; // @[core.scala 24:19]
  wire [31:0] rf_io_rfio_rs_data_bits; // @[core.scala 24:19]
  wire  rf_io_rfio_rt_data_valid; // @[core.scala 24:19]
  wire [31:0] rf_io_rfio_rt_data_bits; // @[core.scala 24:19]
  wire  rf_io_commit_valid; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_pc; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_instr; // @[core.scala 24:19]
  wire  rf_io_commit_ip7; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_0; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_1; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_2; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_3; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_4; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_5; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_6; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_7; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_8; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_9; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_10; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_11; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_12; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_13; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_14; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_15; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_16; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_17; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_18; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_19; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_20; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_21; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_22; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_23; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_24; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_25; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_26; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_27; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_28; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_29; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_30; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_gpr_31; // @[core.scala 24:19]
  wire [4:0] rf_io_commit_rd_idx; // @[core.scala 24:19]
  wire [31:0] rf_io_commit_wdata; // @[core.scala 24:19]
  wire  rf_io_commit_wen; // @[core.scala 24:19]
  wire  rf_io_ex_flush_valid; // @[core.scala 24:19]
  wire  ifu_clock; // @[core.scala 25:19]
  wire  ifu_reset; // @[core.scala 25:19]
  wire  ifu_io_imem_req_ready; // @[core.scala 25:19]
  wire  ifu_io_imem_req_valid; // @[core.scala 25:19]
  wire  ifu_io_imem_req_bits_is_cached; // @[core.scala 25:19]
  wire [31:0] ifu_io_imem_req_bits_addr; // @[core.scala 25:19]
  wire  ifu_io_imem_resp_ready; // @[core.scala 25:19]
  wire  ifu_io_imem_resp_valid; // @[core.scala 25:19]
  wire [31:0] ifu_io_imem_resp_bits_data; // @[core.scala 25:19]
  wire  ifu_io_iaddr_req_ready; // @[core.scala 25:19]
  wire  ifu_io_iaddr_req_valid; // @[core.scala 25:19]
  wire [31:0] ifu_io_iaddr_req_bits_vaddr; // @[core.scala 25:19]
  wire  ifu_io_iaddr_resp_ready; // @[core.scala 25:19]
  wire  ifu_io_iaddr_resp_valid; // @[core.scala 25:19]
  wire [31:0] ifu_io_iaddr_resp_bits_paddr; // @[core.scala 25:19]
  wire  ifu_io_iaddr_resp_bits_is_cached; // @[core.scala 25:19]
  wire [4:0] ifu_io_iaddr_resp_bits_ex_et; // @[core.scala 25:19]
  wire [4:0] ifu_io_iaddr_resp_bits_ex_code; // @[core.scala 25:19]
  wire [31:0] ifu_io_iaddr_resp_bits_ex_addr; // @[core.scala 25:19]
  wire [7:0] ifu_io_iaddr_resp_bits_ex_asid; // @[core.scala 25:19]
  wire  ifu_io_fu_out_ready; // @[core.scala 25:19]
  wire  ifu_io_fu_out_valid; // @[core.scala 25:19]
  wire [31:0] ifu_io_fu_out_bits_pc; // @[core.scala 25:19]
  wire [31:0] ifu_io_fu_out_bits_instr; // @[core.scala 25:19]
  wire [4:0] ifu_io_fu_out_bits_ex_et; // @[core.scala 25:19]
  wire [4:0] ifu_io_fu_out_bits_ex_code; // @[core.scala 25:19]
  wire [31:0] ifu_io_fu_out_bits_ex_addr; // @[core.scala 25:19]
  wire [7:0] ifu_io_fu_out_bits_ex_asid; // @[core.scala 25:19]
  wire  ifu_io_br_flush_valid; // @[core.scala 25:19]
  wire [31:0] ifu_io_br_flush_bits_br_target; // @[core.scala 25:19]
  wire  ifu_io_ex_flush_valid; // @[core.scala 25:19]
  wire [31:0] ifu_io_ex_flush_bits_br_target; // @[core.scala 25:19]
  wire  idu_clock; // @[core.scala 26:19]
  wire  idu_reset; // @[core.scala 26:19]
  wire  idu_io_fu_in_ready; // @[core.scala 26:19]
  wire  idu_io_fu_in_valid; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_in_bits_pc; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_in_bits_instr; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_in_bits_ex_et; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_in_bits_ex_code; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_in_bits_ex_addr; // @[core.scala 26:19]
  wire [7:0] idu_io_fu_in_bits_ex_asid; // @[core.scala 26:19]
  wire  idu_io_fu_out_ready; // @[core.scala 26:19]
  wire  idu_io_fu_out_valid; // @[core.scala 26:19]
  wire  idu_io_fu_out_bits_wb_v; // @[core.scala 26:19]
  wire [7:0] idu_io_fu_out_bits_wb_id; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_out_bits_wb_pc; // @[core.scala 26:19]
  wire [5:0] idu_io_fu_out_bits_wb_instr_op; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_wb_instr_rs_idx; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_wb_instr_rt_idx; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_wb_instr_rd_idx; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_wb_instr_shamt; // @[core.scala 26:19]
  wire [5:0] idu_io_fu_out_bits_wb_instr_func; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_wb_rd_idx; // @[core.scala 26:19]
  wire  idu_io_fu_out_bits_wb_wen; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_out_bits_wb_data; // @[core.scala 26:19]
  wire  idu_io_fu_out_bits_wb_is_ds; // @[core.scala 26:19]
  wire  idu_io_fu_out_bits_wb_is_br; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_out_bits_wb_npc; // @[core.scala 26:19]
  wire [2:0] idu_io_fu_out_bits_ops_fu_type; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_ops_fu_op; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_out_bits_ops_op1; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_out_bits_ops_op2; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_ex_et; // @[core.scala 26:19]
  wire [4:0] idu_io_fu_out_bits_ex_code; // @[core.scala 26:19]
  wire [31:0] idu_io_fu_out_bits_ex_addr; // @[core.scala 26:19]
  wire [7:0] idu_io_fu_out_bits_ex_asid; // @[core.scala 26:19]
  wire  idu_io_br_flush_valid; // @[core.scala 26:19]
  wire [31:0] idu_io_br_flush_bits_br_target; // @[core.scala 26:19]
  wire [4:0] idu_io_rfio_rs_idx; // @[core.scala 26:19]
  wire [4:0] idu_io_rfio_rt_idx; // @[core.scala 26:19]
  wire  idu_io_rfio_wen; // @[core.scala 26:19]
  wire [7:0] idu_io_rfio_wid; // @[core.scala 26:19]
  wire [4:0] idu_io_rfio_rd_idx; // @[core.scala 26:19]
  wire  idu_io_rfio_rs_data_valid; // @[core.scala 26:19]
  wire [31:0] idu_io_rfio_rs_data_bits; // @[core.scala 26:19]
  wire  idu_io_rfio_rt_data_valid; // @[core.scala 26:19]
  wire [31:0] idu_io_rfio_rt_data_bits; // @[core.scala 26:19]
  wire  idu_io_ex_flush_valid; // @[core.scala 26:19]
  wire  exu_clock; // @[core.scala 27:19]
  wire  exu_reset; // @[core.scala 27:19]
  wire  exu_io_fu_in_ready; // @[core.scala 27:19]
  wire  exu_io_fu_in_valid; // @[core.scala 27:19]
  wire  exu_io_fu_in_bits_wb_v; // @[core.scala 27:19]
  wire [7:0] exu_io_fu_in_bits_wb_id; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_in_bits_wb_pc; // @[core.scala 27:19]
  wire [5:0] exu_io_fu_in_bits_wb_instr_op; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_wb_instr_rs_idx; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_wb_instr_rt_idx; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_wb_instr_rd_idx; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_wb_instr_shamt; // @[core.scala 27:19]
  wire [5:0] exu_io_fu_in_bits_wb_instr_func; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_wb_rd_idx; // @[core.scala 27:19]
  wire  exu_io_fu_in_bits_wb_wen; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_in_bits_wb_data; // @[core.scala 27:19]
  wire  exu_io_fu_in_bits_wb_is_ds; // @[core.scala 27:19]
  wire  exu_io_fu_in_bits_wb_is_br; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_in_bits_wb_npc; // @[core.scala 27:19]
  wire [2:0] exu_io_fu_in_bits_ops_fu_type; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_ops_fu_op; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_in_bits_ops_op1; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_in_bits_ops_op2; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_ex_et; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_in_bits_ex_code; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_in_bits_ex_addr; // @[core.scala 27:19]
  wire [7:0] exu_io_fu_in_bits_ex_asid; // @[core.scala 27:19]
  wire  exu_io_fu_out_ready; // @[core.scala 27:19]
  wire  exu_io_fu_out_valid; // @[core.scala 27:19]
  wire  exu_io_fu_out_bits_wb_v; // @[core.scala 27:19]
  wire [7:0] exu_io_fu_out_bits_wb_id; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_out_bits_wb_pc; // @[core.scala 27:19]
  wire [5:0] exu_io_fu_out_bits_wb_instr_op; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_wb_instr_rs_idx; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_wb_instr_rt_idx; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_wb_instr_rd_idx; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_wb_instr_shamt; // @[core.scala 27:19]
  wire [5:0] exu_io_fu_out_bits_wb_instr_func; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_wb_rd_idx; // @[core.scala 27:19]
  wire  exu_io_fu_out_bits_wb_wen; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_out_bits_wb_data; // @[core.scala 27:19]
  wire  exu_io_fu_out_bits_wb_is_ds; // @[core.scala 27:19]
  wire  exu_io_fu_out_bits_wb_is_br; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_out_bits_wb_npc; // @[core.scala 27:19]
  wire [2:0] exu_io_fu_out_bits_ops_fu_type; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_ops_fu_op; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_out_bits_ops_op1; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_out_bits_ops_op2; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_ex_et; // @[core.scala 27:19]
  wire [4:0] exu_io_fu_out_bits_ex_code; // @[core.scala 27:19]
  wire [31:0] exu_io_fu_out_bits_ex_addr; // @[core.scala 27:19]
  wire [7:0] exu_io_fu_out_bits_ex_asid; // @[core.scala 27:19]
  wire [31:0] exu_io_cp0_rport_addr; // @[core.scala 27:19]
  wire [31:0] exu_io_cp0_rport_data; // @[core.scala 27:19]
  wire  exu_io_cp0_wport_valid; // @[core.scala 27:19]
  wire [31:0] exu_io_cp0_wport_bits_addr; // @[core.scala 27:19]
  wire [31:0] exu_io_cp0_wport_bits_data; // @[core.scala 27:19]
  wire [4:0] exu_io_cp0_tlbr_port_index_index; // @[core.scala 27:19]
  wire [15:0] exu_io_cp0_tlbr_port_pagemask_mask; // @[core.scala 27:19]
  wire [18:0] exu_io_cp0_tlbr_port_entry_hi_vpn; // @[core.scala 27:19]
  wire [7:0] exu_io_cp0_tlbr_port_entry_hi_asid; // @[core.scala 27:19]
  wire [19:0] exu_io_cp0_tlbr_port_entry_lo0_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_cp0_tlbr_port_entry_lo0_c; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbr_port_entry_lo0_d; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbr_port_entry_lo0_v; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbr_port_entry_lo0_g; // @[core.scala 27:19]
  wire [19:0] exu_io_cp0_tlbr_port_entry_lo1_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_cp0_tlbr_port_entry_lo1_c; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbr_port_entry_lo1_d; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbr_port_entry_lo1_v; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbr_port_entry_lo1_g; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_valid; // @[core.scala 27:19]
  wire [15:0] exu_io_cp0_tlbw_port_bits_pagemask_mask; // @[core.scala 27:19]
  wire [18:0] exu_io_cp0_tlbw_port_bits_entry_hi_vpn; // @[core.scala 27:19]
  wire [7:0] exu_io_cp0_tlbw_port_bits_entry_hi_asid; // @[core.scala 27:19]
  wire [19:0] exu_io_cp0_tlbw_port_bits_entry_lo0_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_cp0_tlbw_port_bits_entry_lo0_c; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_bits_entry_lo0_d; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_bits_entry_lo0_v; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_bits_entry_lo0_g; // @[core.scala 27:19]
  wire [19:0] exu_io_cp0_tlbw_port_bits_entry_lo1_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_cp0_tlbw_port_bits_entry_lo1_c; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_bits_entry_lo1_d; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_bits_entry_lo1_v; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbw_port_bits_entry_lo1_g; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbp_port_valid; // @[core.scala 27:19]
  wire  exu_io_cp0_tlbp_port_bits_index_p; // @[core.scala 27:19]
  wire [4:0] exu_io_cp0_tlbp_port_bits_index_index; // @[core.scala 27:19]
  wire  exu_io_daddr_req_valid; // @[core.scala 27:19]
  wire  exu_io_daddr_req_bits_func; // @[core.scala 27:19]
  wire [31:0] exu_io_daddr_req_bits_vaddr; // @[core.scala 27:19]
  wire [1:0] exu_io_daddr_req_bits_len; // @[core.scala 27:19]
  wire  exu_io_daddr_req_bits_is_aligned; // @[core.scala 27:19]
  wire [31:0] exu_io_daddr_resp_bits_paddr; // @[core.scala 27:19]
  wire [4:0] exu_io_daddr_resp_bits_ex_et; // @[core.scala 27:19]
  wire [4:0] exu_io_daddr_resp_bits_ex_code; // @[core.scala 27:19]
  wire [31:0] exu_io_daddr_resp_bits_ex_addr; // @[core.scala 27:19]
  wire [7:0] exu_io_daddr_resp_bits_ex_asid; // @[core.scala 27:19]
  wire [4:0] exu_io_tlb_rport_index; // @[core.scala 27:19]
  wire [15:0] exu_io_tlb_rport_entry_pagemask; // @[core.scala 27:19]
  wire [18:0] exu_io_tlb_rport_entry_vpn; // @[core.scala 27:19]
  wire  exu_io_tlb_rport_entry_g; // @[core.scala 27:19]
  wire [7:0] exu_io_tlb_rport_entry_asid; // @[core.scala 27:19]
  wire [23:0] exu_io_tlb_rport_entry_p0_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_tlb_rport_entry_p0_c; // @[core.scala 27:19]
  wire  exu_io_tlb_rport_entry_p0_d; // @[core.scala 27:19]
  wire  exu_io_tlb_rport_entry_p0_v; // @[core.scala 27:19]
  wire [23:0] exu_io_tlb_rport_entry_p1_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_tlb_rport_entry_p1_c; // @[core.scala 27:19]
  wire  exu_io_tlb_rport_entry_p1_d; // @[core.scala 27:19]
  wire  exu_io_tlb_rport_entry_p1_v; // @[core.scala 27:19]
  wire  exu_io_tlb_wport_valid; // @[core.scala 27:19]
  wire [4:0] exu_io_tlb_wport_bits_index; // @[core.scala 27:19]
  wire [15:0] exu_io_tlb_wport_bits_entry_pagemask; // @[core.scala 27:19]
  wire [18:0] exu_io_tlb_wport_bits_entry_vpn; // @[core.scala 27:19]
  wire  exu_io_tlb_wport_bits_entry_g; // @[core.scala 27:19]
  wire [7:0] exu_io_tlb_wport_bits_entry_asid; // @[core.scala 27:19]
  wire [23:0] exu_io_tlb_wport_bits_entry_p0_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_tlb_wport_bits_entry_p0_c; // @[core.scala 27:19]
  wire  exu_io_tlb_wport_bits_entry_p0_d; // @[core.scala 27:19]
  wire  exu_io_tlb_wport_bits_entry_p0_v; // @[core.scala 27:19]
  wire [23:0] exu_io_tlb_wport_bits_entry_p1_pfn; // @[core.scala 27:19]
  wire [2:0] exu_io_tlb_wport_bits_entry_p1_c; // @[core.scala 27:19]
  wire  exu_io_tlb_wport_bits_entry_p1_d; // @[core.scala 27:19]
  wire  exu_io_tlb_wport_bits_entry_p1_v; // @[core.scala 27:19]
  wire [18:0] exu_io_tlb_pport_entry_hi_vpn; // @[core.scala 27:19]
  wire [7:0] exu_io_tlb_pport_entry_hi_asid; // @[core.scala 27:19]
  wire  exu_io_tlb_pport_index_p; // @[core.scala 27:19]
  wire [4:0] exu_io_tlb_pport_index_index; // @[core.scala 27:19]
  wire  exu_io_icache_control_valid; // @[core.scala 27:19]
  wire [2:0] exu_io_icache_control_bits_op; // @[core.scala 27:19]
  wire [31:0] exu_io_icache_control_bits_addr; // @[core.scala 27:19]
  wire  exu_io_bp_valid; // @[core.scala 27:19]
  wire  exu_io_bp_bits_v; // @[core.scala 27:19]
  wire [4:0] exu_io_bp_bits_rd_idx; // @[core.scala 27:19]
  wire  exu_io_bp_bits_wen; // @[core.scala 27:19]
  wire [31:0] exu_io_bp_bits_data; // @[core.scala 27:19]
  wire  exu_io_ex_flush_valid; // @[core.scala 27:19]
  wire  ehu_clock; // @[core.scala 28:19]
  wire  ehu_reset; // @[core.scala 28:19]
  wire  ehu_io_fu_in_ready; // @[core.scala 28:19]
  wire  ehu_io_fu_in_valid; // @[core.scala 28:19]
  wire  ehu_io_fu_in_bits_wb_v; // @[core.scala 28:19]
  wire [7:0] ehu_io_fu_in_bits_wb_id; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_in_bits_wb_pc; // @[core.scala 28:19]
  wire [5:0] ehu_io_fu_in_bits_wb_instr_op; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_wb_instr_rs_idx; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_wb_instr_rt_idx; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_wb_instr_rd_idx; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_wb_instr_shamt; // @[core.scala 28:19]
  wire [5:0] ehu_io_fu_in_bits_wb_instr_func; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_wb_rd_idx; // @[core.scala 28:19]
  wire  ehu_io_fu_in_bits_wb_wen; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_in_bits_wb_data; // @[core.scala 28:19]
  wire  ehu_io_fu_in_bits_wb_is_ds; // @[core.scala 28:19]
  wire  ehu_io_fu_in_bits_wb_is_br; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_in_bits_wb_npc; // @[core.scala 28:19]
  wire [2:0] ehu_io_fu_in_bits_ops_fu_type; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_ops_fu_op; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_in_bits_ops_op1; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_in_bits_ops_op2; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_ex_et; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_in_bits_ex_code; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_in_bits_ex_addr; // @[core.scala 28:19]
  wire [7:0] ehu_io_fu_in_bits_ex_asid; // @[core.scala 28:19]
  wire  ehu_io_fu_out_ready; // @[core.scala 28:19]
  wire  ehu_io_fu_out_valid; // @[core.scala 28:19]
  wire  ehu_io_fu_out_bits_wb_v; // @[core.scala 28:19]
  wire [7:0] ehu_io_fu_out_bits_wb_id; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_out_bits_wb_pc; // @[core.scala 28:19]
  wire [5:0] ehu_io_fu_out_bits_wb_instr_op; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_out_bits_wb_instr_rs_idx; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_out_bits_wb_instr_rt_idx; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_out_bits_wb_instr_rd_idx; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_out_bits_wb_instr_shamt; // @[core.scala 28:19]
  wire [5:0] ehu_io_fu_out_bits_wb_instr_func; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_out_bits_wb_rd_idx; // @[core.scala 28:19]
  wire  ehu_io_fu_out_bits_wb_wen; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_out_bits_wb_data; // @[core.scala 28:19]
  wire  ehu_io_fu_out_bits_wb_ip7; // @[core.scala 28:19]
  wire  ehu_io_fu_out_bits_wb_is_ds; // @[core.scala 28:19]
  wire  ehu_io_fu_out_bits_wb_is_br; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_out_bits_wb_npc; // @[core.scala 28:19]
  wire [2:0] ehu_io_fu_out_bits_ops_fu_type; // @[core.scala 28:19]
  wire [4:0] ehu_io_fu_out_bits_ops_fu_op; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_out_bits_ops_op1; // @[core.scala 28:19]
  wire [31:0] ehu_io_fu_out_bits_ops_op2; // @[core.scala 28:19]
  wire  ehu_io_fu_out_bits_is_cached; // @[core.scala 28:19]
  wire  ehu_io_cp0_valid; // @[core.scala 28:19]
  wire  ehu_io_cp0_ip7; // @[core.scala 28:19]
  wire [4:0] ehu_io_cp0_ex_et; // @[core.scala 28:19]
  wire [4:0] ehu_io_cp0_ex_code; // @[core.scala 28:19]
  wire [31:0] ehu_io_cp0_ex_addr; // @[core.scala 28:19]
  wire [7:0] ehu_io_cp0_ex_asid; // @[core.scala 28:19]
  wire [31:0] ehu_io_cp0_wb_pc; // @[core.scala 28:19]
  wire  ehu_io_cp0_wb_is_ds; // @[core.scala 28:19]
  wire  ehu_io_cp0_wb_is_br; // @[core.scala 28:19]
  wire [31:0] ehu_io_cp0_wb_npc; // @[core.scala 28:19]
  wire  ehu_io_ex_flush_valid; // @[core.scala 28:19]
  wire  cp0_clock; // @[core.scala 29:19]
  wire  cp0_reset; // @[core.scala 29:19]
  wire [31:0] cp0_io_rport_addr; // @[core.scala 29:19]
  wire [31:0] cp0_io_rport_data; // @[core.scala 29:19]
  wire  cp0_io_wport_valid; // @[core.scala 29:19]
  wire [31:0] cp0_io_wport_bits_addr; // @[core.scala 29:19]
  wire [31:0] cp0_io_wport_bits_data; // @[core.scala 29:19]
  wire [4:0] cp0_io_tlbr_port_index_index; // @[core.scala 29:19]
  wire [15:0] cp0_io_tlbr_port_pagemask_mask; // @[core.scala 29:19]
  wire [18:0] cp0_io_tlbr_port_entry_hi_vpn; // @[core.scala 29:19]
  wire [7:0] cp0_io_tlbr_port_entry_hi_asid; // @[core.scala 29:19]
  wire [19:0] cp0_io_tlbr_port_entry_lo0_pfn; // @[core.scala 29:19]
  wire [2:0] cp0_io_tlbr_port_entry_lo0_c; // @[core.scala 29:19]
  wire  cp0_io_tlbr_port_entry_lo0_d; // @[core.scala 29:19]
  wire  cp0_io_tlbr_port_entry_lo0_v; // @[core.scala 29:19]
  wire  cp0_io_tlbr_port_entry_lo0_g; // @[core.scala 29:19]
  wire [19:0] cp0_io_tlbr_port_entry_lo1_pfn; // @[core.scala 29:19]
  wire [2:0] cp0_io_tlbr_port_entry_lo1_c; // @[core.scala 29:19]
  wire  cp0_io_tlbr_port_entry_lo1_d; // @[core.scala 29:19]
  wire  cp0_io_tlbr_port_entry_lo1_v; // @[core.scala 29:19]
  wire  cp0_io_tlbr_port_entry_lo1_g; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_valid; // @[core.scala 29:19]
  wire [15:0] cp0_io_tlbw_port_bits_pagemask_mask; // @[core.scala 29:19]
  wire [18:0] cp0_io_tlbw_port_bits_entry_hi_vpn; // @[core.scala 29:19]
  wire [7:0] cp0_io_tlbw_port_bits_entry_hi_asid; // @[core.scala 29:19]
  wire [19:0] cp0_io_tlbw_port_bits_entry_lo0_pfn; // @[core.scala 29:19]
  wire [2:0] cp0_io_tlbw_port_bits_entry_lo0_c; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_bits_entry_lo0_d; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_bits_entry_lo0_v; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_bits_entry_lo0_g; // @[core.scala 29:19]
  wire [19:0] cp0_io_tlbw_port_bits_entry_lo1_pfn; // @[core.scala 29:19]
  wire [2:0] cp0_io_tlbw_port_bits_entry_lo1_c; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_bits_entry_lo1_d; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_bits_entry_lo1_v; // @[core.scala 29:19]
  wire  cp0_io_tlbw_port_bits_entry_lo1_g; // @[core.scala 29:19]
  wire  cp0_io_tlbp_port_valid; // @[core.scala 29:19]
  wire  cp0_io_tlbp_port_bits_index_p; // @[core.scala 29:19]
  wire [4:0] cp0_io_tlbp_port_bits_index_index; // @[core.scala 29:19]
  wire  cp0_io_status_ERL; // @[core.scala 29:19]
  wire  cp0_io_ehu_valid; // @[core.scala 29:19]
  wire  cp0_io_ehu_ip7; // @[core.scala 29:19]
  wire [4:0] cp0_io_ehu_ex_et; // @[core.scala 29:19]
  wire [4:0] cp0_io_ehu_ex_code; // @[core.scala 29:19]
  wire [31:0] cp0_io_ehu_ex_addr; // @[core.scala 29:19]
  wire [7:0] cp0_io_ehu_ex_asid; // @[core.scala 29:19]
  wire [31:0] cp0_io_ehu_wb_pc; // @[core.scala 29:19]
  wire  cp0_io_ehu_wb_is_ds; // @[core.scala 29:19]
  wire  cp0_io_ehu_wb_is_br; // @[core.scala 29:19]
  wire [31:0] cp0_io_ehu_wb_npc; // @[core.scala 29:19]
  wire  cp0_io_ex_flush_valid; // @[core.scala 29:19]
  wire [31:0] cp0_io_ex_flush_bits_br_target; // @[core.scala 29:19]
  wire  tlb_clock; // @[core.scala 30:19]
  wire  tlb_reset; // @[core.scala 30:19]
  wire  tlb_io_iaddr_req_ready; // @[core.scala 30:19]
  wire  tlb_io_iaddr_req_valid; // @[core.scala 30:19]
  wire [31:0] tlb_io_iaddr_req_bits_vaddr; // @[core.scala 30:19]
  wire  tlb_io_iaddr_resp_ready; // @[core.scala 30:19]
  wire  tlb_io_iaddr_resp_valid; // @[core.scala 30:19]
  wire [31:0] tlb_io_iaddr_resp_bits_paddr; // @[core.scala 30:19]
  wire  tlb_io_iaddr_resp_bits_is_cached; // @[core.scala 30:19]
  wire [4:0] tlb_io_iaddr_resp_bits_ex_et; // @[core.scala 30:19]
  wire [4:0] tlb_io_iaddr_resp_bits_ex_code; // @[core.scala 30:19]
  wire [31:0] tlb_io_iaddr_resp_bits_ex_addr; // @[core.scala 30:19]
  wire [7:0] tlb_io_iaddr_resp_bits_ex_asid; // @[core.scala 30:19]
  wire  tlb_io_daddr_req_ready; // @[core.scala 30:19]
  wire  tlb_io_daddr_req_valid; // @[core.scala 30:19]
  wire  tlb_io_daddr_req_bits_func; // @[core.scala 30:19]
  wire [31:0] tlb_io_daddr_req_bits_vaddr; // @[core.scala 30:19]
  wire [1:0] tlb_io_daddr_req_bits_len; // @[core.scala 30:19]
  wire  tlb_io_daddr_req_bits_is_aligned; // @[core.scala 30:19]
  wire [31:0] tlb_io_daddr_resp_bits_paddr; // @[core.scala 30:19]
  wire [4:0] tlb_io_daddr_resp_bits_ex_et; // @[core.scala 30:19]
  wire [4:0] tlb_io_daddr_resp_bits_ex_code; // @[core.scala 30:19]
  wire [31:0] tlb_io_daddr_resp_bits_ex_addr; // @[core.scala 30:19]
  wire [7:0] tlb_io_daddr_resp_bits_ex_asid; // @[core.scala 30:19]
  wire [4:0] tlb_io_rport_index; // @[core.scala 30:19]
  wire [15:0] tlb_io_rport_entry_pagemask; // @[core.scala 30:19]
  wire [18:0] tlb_io_rport_entry_vpn; // @[core.scala 30:19]
  wire  tlb_io_rport_entry_g; // @[core.scala 30:19]
  wire [7:0] tlb_io_rport_entry_asid; // @[core.scala 30:19]
  wire [23:0] tlb_io_rport_entry_p0_pfn; // @[core.scala 30:19]
  wire [2:0] tlb_io_rport_entry_p0_c; // @[core.scala 30:19]
  wire  tlb_io_rport_entry_p0_d; // @[core.scala 30:19]
  wire  tlb_io_rport_entry_p0_v; // @[core.scala 30:19]
  wire [23:0] tlb_io_rport_entry_p1_pfn; // @[core.scala 30:19]
  wire [2:0] tlb_io_rport_entry_p1_c; // @[core.scala 30:19]
  wire  tlb_io_rport_entry_p1_d; // @[core.scala 30:19]
  wire  tlb_io_rport_entry_p1_v; // @[core.scala 30:19]
  wire  tlb_io_wport_valid; // @[core.scala 30:19]
  wire [4:0] tlb_io_wport_bits_index; // @[core.scala 30:19]
  wire [15:0] tlb_io_wport_bits_entry_pagemask; // @[core.scala 30:19]
  wire [18:0] tlb_io_wport_bits_entry_vpn; // @[core.scala 30:19]
  wire  tlb_io_wport_bits_entry_g; // @[core.scala 30:19]
  wire [7:0] tlb_io_wport_bits_entry_asid; // @[core.scala 30:19]
  wire [23:0] tlb_io_wport_bits_entry_p0_pfn; // @[core.scala 30:19]
  wire [2:0] tlb_io_wport_bits_entry_p0_c; // @[core.scala 30:19]
  wire  tlb_io_wport_bits_entry_p0_d; // @[core.scala 30:19]
  wire  tlb_io_wport_bits_entry_p0_v; // @[core.scala 30:19]
  wire [23:0] tlb_io_wport_bits_entry_p1_pfn; // @[core.scala 30:19]
  wire [2:0] tlb_io_wport_bits_entry_p1_c; // @[core.scala 30:19]
  wire  tlb_io_wport_bits_entry_p1_d; // @[core.scala 30:19]
  wire  tlb_io_wport_bits_entry_p1_v; // @[core.scala 30:19]
  wire [18:0] tlb_io_pport_entry_hi_vpn; // @[core.scala 30:19]
  wire [7:0] tlb_io_pport_entry_hi_asid; // @[core.scala 30:19]
  wire  tlb_io_pport_index_p; // @[core.scala 30:19]
  wire [4:0] tlb_io_pport_index_index; // @[core.scala 30:19]
  wire  tlb_io_status_ERL; // @[core.scala 30:19]
  wire  tlb_io_br_flush_valid; // @[core.scala 30:19]
  wire  tlb_io_ex_flush_valid; // @[core.scala 30:19]
  wire  msu_clock; // @[core.scala 31:19]
  wire  msu_reset; // @[core.scala 31:19]
  wire  msu_io_fu_in_ready; // @[core.scala 31:19]
  wire  msu_io_fu_in_valid; // @[core.scala 31:19]
  wire  msu_io_fu_in_bits_wb_v; // @[core.scala 31:19]
  wire [7:0] msu_io_fu_in_bits_wb_id; // @[core.scala 31:19]
  wire [31:0] msu_io_fu_in_bits_wb_pc; // @[core.scala 31:19]
  wire [5:0] msu_io_fu_in_bits_wb_instr_op; // @[core.scala 31:19]
  wire [4:0] msu_io_fu_in_bits_wb_instr_rs_idx; // @[core.scala 31:19]
  wire [4:0] msu_io_fu_in_bits_wb_instr_rt_idx; // @[core.scala 31:19]
  wire [4:0] msu_io_fu_in_bits_wb_instr_rd_idx; // @[core.scala 31:19]
  wire [4:0] msu_io_fu_in_bits_wb_instr_shamt; // @[core.scala 31:19]
  wire [5:0] msu_io_fu_in_bits_wb_instr_func; // @[core.scala 31:19]
  wire [4:0] msu_io_fu_in_bits_wb_rd_idx; // @[core.scala 31:19]
  wire  msu_io_fu_in_bits_wb_wen; // @[core.scala 31:19]
  wire [31:0] msu_io_fu_in_bits_wb_data; // @[core.scala 31:19]
  wire  msu_io_fu_in_bits_wb_ip7; // @[core.scala 31:19]
  wire  msu_io_fu_in_bits_wb_is_ds; // @[core.scala 31:19]
  wire  msu_io_fu_in_bits_wb_is_br; // @[core.scala 31:19]
  wire [31:0] msu_io_fu_in_bits_wb_npc; // @[core.scala 31:19]
  wire [2:0] msu_io_fu_in_bits_ops_fu_type; // @[core.scala 31:19]
  wire [4:0] msu_io_fu_in_bits_ops_fu_op; // @[core.scala 31:19]
  wire [31:0] msu_io_fu_in_bits_ops_op1; // @[core.scala 31:19]
  wire [31:0] msu_io_fu_in_bits_ops_op2; // @[core.scala 31:19]
  wire  msu_io_fu_in_bits_is_cached; // @[core.scala 31:19]
  wire  msu_io_wb_valid; // @[core.scala 31:19]
  wire  msu_io_wb_bits_v; // @[core.scala 31:19]
  wire [7:0] msu_io_wb_bits_id; // @[core.scala 31:19]
  wire [31:0] msu_io_wb_bits_pc; // @[core.scala 31:19]
  wire [5:0] msu_io_wb_bits_instr_op; // @[core.scala 31:19]
  wire [4:0] msu_io_wb_bits_instr_rs_idx; // @[core.scala 31:19]
  wire [4:0] msu_io_wb_bits_instr_rt_idx; // @[core.scala 31:19]
  wire [4:0] msu_io_wb_bits_instr_rd_idx; // @[core.scala 31:19]
  wire [4:0] msu_io_wb_bits_instr_shamt; // @[core.scala 31:19]
  wire [5:0] msu_io_wb_bits_instr_func; // @[core.scala 31:19]
  wire [4:0] msu_io_wb_bits_rd_idx; // @[core.scala 31:19]
  wire  msu_io_wb_bits_wen; // @[core.scala 31:19]
  wire [31:0] msu_io_wb_bits_data; // @[core.scala 31:19]
  wire  msu_io_wb_bits_ip7; // @[core.scala 31:19]
  wire  msu_io_divider_data_dividend_tvalid; // @[core.scala 31:19]
  wire  msu_io_divider_data_divisor_tvalid; // @[core.scala 31:19]
  wire  msu_io_divider_data_dout_tvalid; // @[core.scala 31:19]
  wire [39:0] msu_io_divider_data_dividend_tdata; // @[core.scala 31:19]
  wire [39:0] msu_io_divider_data_divisor_tdata; // @[core.scala 31:19]
  wire [79:0] msu_io_divider_data_dout_tdata; // @[core.scala 31:19]
  wire [32:0] msu_io_multiplier_data_a; // @[core.scala 31:19]
  wire [32:0] msu_io_multiplier_data_b; // @[core.scala 31:19]
  wire [65:0] msu_io_multiplier_data_dout; // @[core.scala 31:19]
  wire  msu_io_dmem_req_ready; // @[core.scala 31:19]
  wire  msu_io_dmem_req_valid; // @[core.scala 31:19]
  wire  msu_io_dmem_req_bits_is_cached; // @[core.scala 31:19]
  wire [31:0] msu_io_dmem_req_bits_addr; // @[core.scala 31:19]
  wire [1:0] msu_io_dmem_req_bits_len; // @[core.scala 31:19]
  wire [3:0] msu_io_dmem_req_bits_strb; // @[core.scala 31:19]
  wire [31:0] msu_io_dmem_req_bits_data; // @[core.scala 31:19]
  wire  msu_io_dmem_req_bits_func; // @[core.scala 31:19]
  wire  msu_io_dmem_resp_valid; // @[core.scala 31:19]
  wire [31:0] msu_io_dmem_resp_bits_data; // @[core.scala 31:19]
  RegFile rf ( // @[core.scala 24:19]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_bp_valid(rf_io_bp_valid),
    .io_bp_bits_v(rf_io_bp_bits_v),
    .io_bp_bits_rd_idx(rf_io_bp_bits_rd_idx),
    .io_bp_bits_wen(rf_io_bp_bits_wen),
    .io_bp_bits_data(rf_io_bp_bits_data),
    .io_wb_valid(rf_io_wb_valid),
    .io_wb_bits_v(rf_io_wb_bits_v),
    .io_wb_bits_id(rf_io_wb_bits_id),
    .io_wb_bits_pc(rf_io_wb_bits_pc),
    .io_wb_bits_instr_op(rf_io_wb_bits_instr_op),
    .io_wb_bits_instr_rs_idx(rf_io_wb_bits_instr_rs_idx),
    .io_wb_bits_instr_rt_idx(rf_io_wb_bits_instr_rt_idx),
    .io_wb_bits_instr_rd_idx(rf_io_wb_bits_instr_rd_idx),
    .io_wb_bits_instr_shamt(rf_io_wb_bits_instr_shamt),
    .io_wb_bits_instr_func(rf_io_wb_bits_instr_func),
    .io_wb_bits_rd_idx(rf_io_wb_bits_rd_idx),
    .io_wb_bits_wen(rf_io_wb_bits_wen),
    .io_wb_bits_data(rf_io_wb_bits_data),
    .io_wb_bits_ip7(rf_io_wb_bits_ip7),
    .io_rfio_rs_idx(rf_io_rfio_rs_idx),
    .io_rfio_rt_idx(rf_io_rfio_rt_idx),
    .io_rfio_wen(rf_io_rfio_wen),
    .io_rfio_wid(rf_io_rfio_wid),
    .io_rfio_rd_idx(rf_io_rfio_rd_idx),
    .io_rfio_rs_data_valid(rf_io_rfio_rs_data_valid),
    .io_rfio_rs_data_bits(rf_io_rfio_rs_data_bits),
    .io_rfio_rt_data_valid(rf_io_rfio_rt_data_valid),
    .io_rfio_rt_data_bits(rf_io_rfio_rt_data_bits),
    .io_commit_valid(rf_io_commit_valid),
    .io_commit_pc(rf_io_commit_pc),
    .io_commit_instr(rf_io_commit_instr),
    .io_commit_ip7(rf_io_commit_ip7),
    .io_commit_gpr_0(rf_io_commit_gpr_0),
    .io_commit_gpr_1(rf_io_commit_gpr_1),
    .io_commit_gpr_2(rf_io_commit_gpr_2),
    .io_commit_gpr_3(rf_io_commit_gpr_3),
    .io_commit_gpr_4(rf_io_commit_gpr_4),
    .io_commit_gpr_5(rf_io_commit_gpr_5),
    .io_commit_gpr_6(rf_io_commit_gpr_6),
    .io_commit_gpr_7(rf_io_commit_gpr_7),
    .io_commit_gpr_8(rf_io_commit_gpr_8),
    .io_commit_gpr_9(rf_io_commit_gpr_9),
    .io_commit_gpr_10(rf_io_commit_gpr_10),
    .io_commit_gpr_11(rf_io_commit_gpr_11),
    .io_commit_gpr_12(rf_io_commit_gpr_12),
    .io_commit_gpr_13(rf_io_commit_gpr_13),
    .io_commit_gpr_14(rf_io_commit_gpr_14),
    .io_commit_gpr_15(rf_io_commit_gpr_15),
    .io_commit_gpr_16(rf_io_commit_gpr_16),
    .io_commit_gpr_17(rf_io_commit_gpr_17),
    .io_commit_gpr_18(rf_io_commit_gpr_18),
    .io_commit_gpr_19(rf_io_commit_gpr_19),
    .io_commit_gpr_20(rf_io_commit_gpr_20),
    .io_commit_gpr_21(rf_io_commit_gpr_21),
    .io_commit_gpr_22(rf_io_commit_gpr_22),
    .io_commit_gpr_23(rf_io_commit_gpr_23),
    .io_commit_gpr_24(rf_io_commit_gpr_24),
    .io_commit_gpr_25(rf_io_commit_gpr_25),
    .io_commit_gpr_26(rf_io_commit_gpr_26),
    .io_commit_gpr_27(rf_io_commit_gpr_27),
    .io_commit_gpr_28(rf_io_commit_gpr_28),
    .io_commit_gpr_29(rf_io_commit_gpr_29),
    .io_commit_gpr_30(rf_io_commit_gpr_30),
    .io_commit_gpr_31(rf_io_commit_gpr_31),
    .io_commit_rd_idx(rf_io_commit_rd_idx),
    .io_commit_wdata(rf_io_commit_wdata),
    .io_commit_wen(rf_io_commit_wen),
    .io_ex_flush_valid(rf_io_ex_flush_valid)
  );
  IFU ifu ( // @[core.scala 25:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_is_cached(ifu_io_imem_req_bits_is_cached),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_data(ifu_io_imem_resp_bits_data),
    .io_iaddr_req_ready(ifu_io_iaddr_req_ready),
    .io_iaddr_req_valid(ifu_io_iaddr_req_valid),
    .io_iaddr_req_bits_vaddr(ifu_io_iaddr_req_bits_vaddr),
    .io_iaddr_resp_ready(ifu_io_iaddr_resp_ready),
    .io_iaddr_resp_valid(ifu_io_iaddr_resp_valid),
    .io_iaddr_resp_bits_paddr(ifu_io_iaddr_resp_bits_paddr),
    .io_iaddr_resp_bits_is_cached(ifu_io_iaddr_resp_bits_is_cached),
    .io_iaddr_resp_bits_ex_et(ifu_io_iaddr_resp_bits_ex_et),
    .io_iaddr_resp_bits_ex_code(ifu_io_iaddr_resp_bits_ex_code),
    .io_iaddr_resp_bits_ex_addr(ifu_io_iaddr_resp_bits_ex_addr),
    .io_iaddr_resp_bits_ex_asid(ifu_io_iaddr_resp_bits_ex_asid),
    .io_fu_out_ready(ifu_io_fu_out_ready),
    .io_fu_out_valid(ifu_io_fu_out_valid),
    .io_fu_out_bits_pc(ifu_io_fu_out_bits_pc),
    .io_fu_out_bits_instr(ifu_io_fu_out_bits_instr),
    .io_fu_out_bits_ex_et(ifu_io_fu_out_bits_ex_et),
    .io_fu_out_bits_ex_code(ifu_io_fu_out_bits_ex_code),
    .io_fu_out_bits_ex_addr(ifu_io_fu_out_bits_ex_addr),
    .io_fu_out_bits_ex_asid(ifu_io_fu_out_bits_ex_asid),
    .io_br_flush_valid(ifu_io_br_flush_valid),
    .io_br_flush_bits_br_target(ifu_io_br_flush_bits_br_target),
    .io_ex_flush_valid(ifu_io_ex_flush_valid),
    .io_ex_flush_bits_br_target(ifu_io_ex_flush_bits_br_target)
  );
  IDU idu ( // @[core.scala 26:19]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_fu_in_ready(idu_io_fu_in_ready),
    .io_fu_in_valid(idu_io_fu_in_valid),
    .io_fu_in_bits_pc(idu_io_fu_in_bits_pc),
    .io_fu_in_bits_instr(idu_io_fu_in_bits_instr),
    .io_fu_in_bits_ex_et(idu_io_fu_in_bits_ex_et),
    .io_fu_in_bits_ex_code(idu_io_fu_in_bits_ex_code),
    .io_fu_in_bits_ex_addr(idu_io_fu_in_bits_ex_addr),
    .io_fu_in_bits_ex_asid(idu_io_fu_in_bits_ex_asid),
    .io_fu_out_ready(idu_io_fu_out_ready),
    .io_fu_out_valid(idu_io_fu_out_valid),
    .io_fu_out_bits_wb_v(idu_io_fu_out_bits_wb_v),
    .io_fu_out_bits_wb_id(idu_io_fu_out_bits_wb_id),
    .io_fu_out_bits_wb_pc(idu_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(idu_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(idu_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(idu_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(idu_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(idu_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(idu_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_rd_idx(idu_io_fu_out_bits_wb_rd_idx),
    .io_fu_out_bits_wb_wen(idu_io_fu_out_bits_wb_wen),
    .io_fu_out_bits_wb_data(idu_io_fu_out_bits_wb_data),
    .io_fu_out_bits_wb_is_ds(idu_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_wb_is_br(idu_io_fu_out_bits_wb_is_br),
    .io_fu_out_bits_wb_npc(idu_io_fu_out_bits_wb_npc),
    .io_fu_out_bits_ops_fu_type(idu_io_fu_out_bits_ops_fu_type),
    .io_fu_out_bits_ops_fu_op(idu_io_fu_out_bits_ops_fu_op),
    .io_fu_out_bits_ops_op1(idu_io_fu_out_bits_ops_op1),
    .io_fu_out_bits_ops_op2(idu_io_fu_out_bits_ops_op2),
    .io_fu_out_bits_ex_et(idu_io_fu_out_bits_ex_et),
    .io_fu_out_bits_ex_code(idu_io_fu_out_bits_ex_code),
    .io_fu_out_bits_ex_addr(idu_io_fu_out_bits_ex_addr),
    .io_fu_out_bits_ex_asid(idu_io_fu_out_bits_ex_asid),
    .io_br_flush_valid(idu_io_br_flush_valid),
    .io_br_flush_bits_br_target(idu_io_br_flush_bits_br_target),
    .io_rfio_rs_idx(idu_io_rfio_rs_idx),
    .io_rfio_rt_idx(idu_io_rfio_rt_idx),
    .io_rfio_wen(idu_io_rfio_wen),
    .io_rfio_wid(idu_io_rfio_wid),
    .io_rfio_rd_idx(idu_io_rfio_rd_idx),
    .io_rfio_rs_data_valid(idu_io_rfio_rs_data_valid),
    .io_rfio_rs_data_bits(idu_io_rfio_rs_data_bits),
    .io_rfio_rt_data_valid(idu_io_rfio_rt_data_valid),
    .io_rfio_rt_data_bits(idu_io_rfio_rt_data_bits),
    .io_ex_flush_valid(idu_io_ex_flush_valid)
  );
  EXU exu ( // @[core.scala 27:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_fu_in_ready(exu_io_fu_in_ready),
    .io_fu_in_valid(exu_io_fu_in_valid),
    .io_fu_in_bits_wb_v(exu_io_fu_in_bits_wb_v),
    .io_fu_in_bits_wb_id(exu_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(exu_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(exu_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(exu_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(exu_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(exu_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(exu_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(exu_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(exu_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_wen(exu_io_fu_in_bits_wb_wen),
    .io_fu_in_bits_wb_data(exu_io_fu_in_bits_wb_data),
    .io_fu_in_bits_wb_is_ds(exu_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(exu_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(exu_io_fu_in_bits_wb_npc),
    .io_fu_in_bits_ops_fu_type(exu_io_fu_in_bits_ops_fu_type),
    .io_fu_in_bits_ops_fu_op(exu_io_fu_in_bits_ops_fu_op),
    .io_fu_in_bits_ops_op1(exu_io_fu_in_bits_ops_op1),
    .io_fu_in_bits_ops_op2(exu_io_fu_in_bits_ops_op2),
    .io_fu_in_bits_ex_et(exu_io_fu_in_bits_ex_et),
    .io_fu_in_bits_ex_code(exu_io_fu_in_bits_ex_code),
    .io_fu_in_bits_ex_addr(exu_io_fu_in_bits_ex_addr),
    .io_fu_in_bits_ex_asid(exu_io_fu_in_bits_ex_asid),
    .io_fu_out_ready(exu_io_fu_out_ready),
    .io_fu_out_valid(exu_io_fu_out_valid),
    .io_fu_out_bits_wb_v(exu_io_fu_out_bits_wb_v),
    .io_fu_out_bits_wb_id(exu_io_fu_out_bits_wb_id),
    .io_fu_out_bits_wb_pc(exu_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(exu_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(exu_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(exu_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(exu_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(exu_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(exu_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_rd_idx(exu_io_fu_out_bits_wb_rd_idx),
    .io_fu_out_bits_wb_wen(exu_io_fu_out_bits_wb_wen),
    .io_fu_out_bits_wb_data(exu_io_fu_out_bits_wb_data),
    .io_fu_out_bits_wb_is_ds(exu_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_wb_is_br(exu_io_fu_out_bits_wb_is_br),
    .io_fu_out_bits_wb_npc(exu_io_fu_out_bits_wb_npc),
    .io_fu_out_bits_ops_fu_type(exu_io_fu_out_bits_ops_fu_type),
    .io_fu_out_bits_ops_fu_op(exu_io_fu_out_bits_ops_fu_op),
    .io_fu_out_bits_ops_op1(exu_io_fu_out_bits_ops_op1),
    .io_fu_out_bits_ops_op2(exu_io_fu_out_bits_ops_op2),
    .io_fu_out_bits_ex_et(exu_io_fu_out_bits_ex_et),
    .io_fu_out_bits_ex_code(exu_io_fu_out_bits_ex_code),
    .io_fu_out_bits_ex_addr(exu_io_fu_out_bits_ex_addr),
    .io_fu_out_bits_ex_asid(exu_io_fu_out_bits_ex_asid),
    .io_cp0_rport_addr(exu_io_cp0_rport_addr),
    .io_cp0_rport_data(exu_io_cp0_rport_data),
    .io_cp0_wport_valid(exu_io_cp0_wport_valid),
    .io_cp0_wport_bits_addr(exu_io_cp0_wport_bits_addr),
    .io_cp0_wport_bits_data(exu_io_cp0_wport_bits_data),
    .io_cp0_tlbr_port_index_index(exu_io_cp0_tlbr_port_index_index),
    .io_cp0_tlbr_port_pagemask_mask(exu_io_cp0_tlbr_port_pagemask_mask),
    .io_cp0_tlbr_port_entry_hi_vpn(exu_io_cp0_tlbr_port_entry_hi_vpn),
    .io_cp0_tlbr_port_entry_hi_asid(exu_io_cp0_tlbr_port_entry_hi_asid),
    .io_cp0_tlbr_port_entry_lo0_pfn(exu_io_cp0_tlbr_port_entry_lo0_pfn),
    .io_cp0_tlbr_port_entry_lo0_c(exu_io_cp0_tlbr_port_entry_lo0_c),
    .io_cp0_tlbr_port_entry_lo0_d(exu_io_cp0_tlbr_port_entry_lo0_d),
    .io_cp0_tlbr_port_entry_lo0_v(exu_io_cp0_tlbr_port_entry_lo0_v),
    .io_cp0_tlbr_port_entry_lo0_g(exu_io_cp0_tlbr_port_entry_lo0_g),
    .io_cp0_tlbr_port_entry_lo1_pfn(exu_io_cp0_tlbr_port_entry_lo1_pfn),
    .io_cp0_tlbr_port_entry_lo1_c(exu_io_cp0_tlbr_port_entry_lo1_c),
    .io_cp0_tlbr_port_entry_lo1_d(exu_io_cp0_tlbr_port_entry_lo1_d),
    .io_cp0_tlbr_port_entry_lo1_v(exu_io_cp0_tlbr_port_entry_lo1_v),
    .io_cp0_tlbr_port_entry_lo1_g(exu_io_cp0_tlbr_port_entry_lo1_g),
    .io_cp0_tlbw_port_valid(exu_io_cp0_tlbw_port_valid),
    .io_cp0_tlbw_port_bits_pagemask_mask(exu_io_cp0_tlbw_port_bits_pagemask_mask),
    .io_cp0_tlbw_port_bits_entry_hi_vpn(exu_io_cp0_tlbw_port_bits_entry_hi_vpn),
    .io_cp0_tlbw_port_bits_entry_hi_asid(exu_io_cp0_tlbw_port_bits_entry_hi_asid),
    .io_cp0_tlbw_port_bits_entry_lo0_pfn(exu_io_cp0_tlbw_port_bits_entry_lo0_pfn),
    .io_cp0_tlbw_port_bits_entry_lo0_c(exu_io_cp0_tlbw_port_bits_entry_lo0_c),
    .io_cp0_tlbw_port_bits_entry_lo0_d(exu_io_cp0_tlbw_port_bits_entry_lo0_d),
    .io_cp0_tlbw_port_bits_entry_lo0_v(exu_io_cp0_tlbw_port_bits_entry_lo0_v),
    .io_cp0_tlbw_port_bits_entry_lo0_g(exu_io_cp0_tlbw_port_bits_entry_lo0_g),
    .io_cp0_tlbw_port_bits_entry_lo1_pfn(exu_io_cp0_tlbw_port_bits_entry_lo1_pfn),
    .io_cp0_tlbw_port_bits_entry_lo1_c(exu_io_cp0_tlbw_port_bits_entry_lo1_c),
    .io_cp0_tlbw_port_bits_entry_lo1_d(exu_io_cp0_tlbw_port_bits_entry_lo1_d),
    .io_cp0_tlbw_port_bits_entry_lo1_v(exu_io_cp0_tlbw_port_bits_entry_lo1_v),
    .io_cp0_tlbw_port_bits_entry_lo1_g(exu_io_cp0_tlbw_port_bits_entry_lo1_g),
    .io_cp0_tlbp_port_valid(exu_io_cp0_tlbp_port_valid),
    .io_cp0_tlbp_port_bits_index_p(exu_io_cp0_tlbp_port_bits_index_p),
    .io_cp0_tlbp_port_bits_index_index(exu_io_cp0_tlbp_port_bits_index_index),
    .io_daddr_req_valid(exu_io_daddr_req_valid),
    .io_daddr_req_bits_func(exu_io_daddr_req_bits_func),
    .io_daddr_req_bits_vaddr(exu_io_daddr_req_bits_vaddr),
    .io_daddr_req_bits_len(exu_io_daddr_req_bits_len),
    .io_daddr_req_bits_is_aligned(exu_io_daddr_req_bits_is_aligned),
    .io_daddr_resp_bits_paddr(exu_io_daddr_resp_bits_paddr),
    .io_daddr_resp_bits_ex_et(exu_io_daddr_resp_bits_ex_et),
    .io_daddr_resp_bits_ex_code(exu_io_daddr_resp_bits_ex_code),
    .io_daddr_resp_bits_ex_addr(exu_io_daddr_resp_bits_ex_addr),
    .io_daddr_resp_bits_ex_asid(exu_io_daddr_resp_bits_ex_asid),
    .io_tlb_rport_index(exu_io_tlb_rport_index),
    .io_tlb_rport_entry_pagemask(exu_io_tlb_rport_entry_pagemask),
    .io_tlb_rport_entry_vpn(exu_io_tlb_rport_entry_vpn),
    .io_tlb_rport_entry_g(exu_io_tlb_rport_entry_g),
    .io_tlb_rport_entry_asid(exu_io_tlb_rport_entry_asid),
    .io_tlb_rport_entry_p0_pfn(exu_io_tlb_rport_entry_p0_pfn),
    .io_tlb_rport_entry_p0_c(exu_io_tlb_rport_entry_p0_c),
    .io_tlb_rport_entry_p0_d(exu_io_tlb_rport_entry_p0_d),
    .io_tlb_rport_entry_p0_v(exu_io_tlb_rport_entry_p0_v),
    .io_tlb_rport_entry_p1_pfn(exu_io_tlb_rport_entry_p1_pfn),
    .io_tlb_rport_entry_p1_c(exu_io_tlb_rport_entry_p1_c),
    .io_tlb_rport_entry_p1_d(exu_io_tlb_rport_entry_p1_d),
    .io_tlb_rport_entry_p1_v(exu_io_tlb_rport_entry_p1_v),
    .io_tlb_wport_valid(exu_io_tlb_wport_valid),
    .io_tlb_wport_bits_index(exu_io_tlb_wport_bits_index),
    .io_tlb_wport_bits_entry_pagemask(exu_io_tlb_wport_bits_entry_pagemask),
    .io_tlb_wport_bits_entry_vpn(exu_io_tlb_wport_bits_entry_vpn),
    .io_tlb_wport_bits_entry_g(exu_io_tlb_wport_bits_entry_g),
    .io_tlb_wport_bits_entry_asid(exu_io_tlb_wport_bits_entry_asid),
    .io_tlb_wport_bits_entry_p0_pfn(exu_io_tlb_wport_bits_entry_p0_pfn),
    .io_tlb_wport_bits_entry_p0_c(exu_io_tlb_wport_bits_entry_p0_c),
    .io_tlb_wport_bits_entry_p0_d(exu_io_tlb_wport_bits_entry_p0_d),
    .io_tlb_wport_bits_entry_p0_v(exu_io_tlb_wport_bits_entry_p0_v),
    .io_tlb_wport_bits_entry_p1_pfn(exu_io_tlb_wport_bits_entry_p1_pfn),
    .io_tlb_wport_bits_entry_p1_c(exu_io_tlb_wport_bits_entry_p1_c),
    .io_tlb_wport_bits_entry_p1_d(exu_io_tlb_wport_bits_entry_p1_d),
    .io_tlb_wport_bits_entry_p1_v(exu_io_tlb_wport_bits_entry_p1_v),
    .io_tlb_pport_entry_hi_vpn(exu_io_tlb_pport_entry_hi_vpn),
    .io_tlb_pport_entry_hi_asid(exu_io_tlb_pport_entry_hi_asid),
    .io_tlb_pport_index_p(exu_io_tlb_pport_index_p),
    .io_tlb_pport_index_index(exu_io_tlb_pport_index_index),
    .io_icache_control_valid(exu_io_icache_control_valid),
    .io_icache_control_bits_op(exu_io_icache_control_bits_op),
    .io_icache_control_bits_addr(exu_io_icache_control_bits_addr),
    .io_bp_valid(exu_io_bp_valid),
    .io_bp_bits_v(exu_io_bp_bits_v),
    .io_bp_bits_rd_idx(exu_io_bp_bits_rd_idx),
    .io_bp_bits_wen(exu_io_bp_bits_wen),
    .io_bp_bits_data(exu_io_bp_bits_data),
    .io_ex_flush_valid(exu_io_ex_flush_valid)
  );
  EHU ehu ( // @[core.scala 28:19]
    .clock(ehu_clock),
    .reset(ehu_reset),
    .io_fu_in_ready(ehu_io_fu_in_ready),
    .io_fu_in_valid(ehu_io_fu_in_valid),
    .io_fu_in_bits_wb_v(ehu_io_fu_in_bits_wb_v),
    .io_fu_in_bits_wb_id(ehu_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(ehu_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(ehu_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(ehu_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(ehu_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(ehu_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(ehu_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(ehu_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(ehu_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_wen(ehu_io_fu_in_bits_wb_wen),
    .io_fu_in_bits_wb_data(ehu_io_fu_in_bits_wb_data),
    .io_fu_in_bits_wb_is_ds(ehu_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(ehu_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(ehu_io_fu_in_bits_wb_npc),
    .io_fu_in_bits_ops_fu_type(ehu_io_fu_in_bits_ops_fu_type),
    .io_fu_in_bits_ops_fu_op(ehu_io_fu_in_bits_ops_fu_op),
    .io_fu_in_bits_ops_op1(ehu_io_fu_in_bits_ops_op1),
    .io_fu_in_bits_ops_op2(ehu_io_fu_in_bits_ops_op2),
    .io_fu_in_bits_ex_et(ehu_io_fu_in_bits_ex_et),
    .io_fu_in_bits_ex_code(ehu_io_fu_in_bits_ex_code),
    .io_fu_in_bits_ex_addr(ehu_io_fu_in_bits_ex_addr),
    .io_fu_in_bits_ex_asid(ehu_io_fu_in_bits_ex_asid),
    .io_fu_out_ready(ehu_io_fu_out_ready),
    .io_fu_out_valid(ehu_io_fu_out_valid),
    .io_fu_out_bits_wb_v(ehu_io_fu_out_bits_wb_v),
    .io_fu_out_bits_wb_id(ehu_io_fu_out_bits_wb_id),
    .io_fu_out_bits_wb_pc(ehu_io_fu_out_bits_wb_pc),
    .io_fu_out_bits_wb_instr_op(ehu_io_fu_out_bits_wb_instr_op),
    .io_fu_out_bits_wb_instr_rs_idx(ehu_io_fu_out_bits_wb_instr_rs_idx),
    .io_fu_out_bits_wb_instr_rt_idx(ehu_io_fu_out_bits_wb_instr_rt_idx),
    .io_fu_out_bits_wb_instr_rd_idx(ehu_io_fu_out_bits_wb_instr_rd_idx),
    .io_fu_out_bits_wb_instr_shamt(ehu_io_fu_out_bits_wb_instr_shamt),
    .io_fu_out_bits_wb_instr_func(ehu_io_fu_out_bits_wb_instr_func),
    .io_fu_out_bits_wb_rd_idx(ehu_io_fu_out_bits_wb_rd_idx),
    .io_fu_out_bits_wb_wen(ehu_io_fu_out_bits_wb_wen),
    .io_fu_out_bits_wb_data(ehu_io_fu_out_bits_wb_data),
    .io_fu_out_bits_wb_ip7(ehu_io_fu_out_bits_wb_ip7),
    .io_fu_out_bits_wb_is_ds(ehu_io_fu_out_bits_wb_is_ds),
    .io_fu_out_bits_wb_is_br(ehu_io_fu_out_bits_wb_is_br),
    .io_fu_out_bits_wb_npc(ehu_io_fu_out_bits_wb_npc),
    .io_fu_out_bits_ops_fu_type(ehu_io_fu_out_bits_ops_fu_type),
    .io_fu_out_bits_ops_fu_op(ehu_io_fu_out_bits_ops_fu_op),
    .io_fu_out_bits_ops_op1(ehu_io_fu_out_bits_ops_op1),
    .io_fu_out_bits_ops_op2(ehu_io_fu_out_bits_ops_op2),
    .io_fu_out_bits_is_cached(ehu_io_fu_out_bits_is_cached),
    .io_cp0_valid(ehu_io_cp0_valid),
    .io_cp0_ip7(ehu_io_cp0_ip7),
    .io_cp0_ex_et(ehu_io_cp0_ex_et),
    .io_cp0_ex_code(ehu_io_cp0_ex_code),
    .io_cp0_ex_addr(ehu_io_cp0_ex_addr),
    .io_cp0_ex_asid(ehu_io_cp0_ex_asid),
    .io_cp0_wb_pc(ehu_io_cp0_wb_pc),
    .io_cp0_wb_is_ds(ehu_io_cp0_wb_is_ds),
    .io_cp0_wb_is_br(ehu_io_cp0_wb_is_br),
    .io_cp0_wb_npc(ehu_io_cp0_wb_npc),
    .io_ex_flush_valid(ehu_io_ex_flush_valid)
  );
  CP0 cp0 ( // @[core.scala 29:19]
    .clock(cp0_clock),
    .reset(cp0_reset),
    .io_rport_addr(cp0_io_rport_addr),
    .io_rport_data(cp0_io_rport_data),
    .io_wport_valid(cp0_io_wport_valid),
    .io_wport_bits_addr(cp0_io_wport_bits_addr),
    .io_wport_bits_data(cp0_io_wport_bits_data),
    .io_tlbr_port_index_index(cp0_io_tlbr_port_index_index),
    .io_tlbr_port_pagemask_mask(cp0_io_tlbr_port_pagemask_mask),
    .io_tlbr_port_entry_hi_vpn(cp0_io_tlbr_port_entry_hi_vpn),
    .io_tlbr_port_entry_hi_asid(cp0_io_tlbr_port_entry_hi_asid),
    .io_tlbr_port_entry_lo0_pfn(cp0_io_tlbr_port_entry_lo0_pfn),
    .io_tlbr_port_entry_lo0_c(cp0_io_tlbr_port_entry_lo0_c),
    .io_tlbr_port_entry_lo0_d(cp0_io_tlbr_port_entry_lo0_d),
    .io_tlbr_port_entry_lo0_v(cp0_io_tlbr_port_entry_lo0_v),
    .io_tlbr_port_entry_lo0_g(cp0_io_tlbr_port_entry_lo0_g),
    .io_tlbr_port_entry_lo1_pfn(cp0_io_tlbr_port_entry_lo1_pfn),
    .io_tlbr_port_entry_lo1_c(cp0_io_tlbr_port_entry_lo1_c),
    .io_tlbr_port_entry_lo1_d(cp0_io_tlbr_port_entry_lo1_d),
    .io_tlbr_port_entry_lo1_v(cp0_io_tlbr_port_entry_lo1_v),
    .io_tlbr_port_entry_lo1_g(cp0_io_tlbr_port_entry_lo1_g),
    .io_tlbw_port_valid(cp0_io_tlbw_port_valid),
    .io_tlbw_port_bits_pagemask_mask(cp0_io_tlbw_port_bits_pagemask_mask),
    .io_tlbw_port_bits_entry_hi_vpn(cp0_io_tlbw_port_bits_entry_hi_vpn),
    .io_tlbw_port_bits_entry_hi_asid(cp0_io_tlbw_port_bits_entry_hi_asid),
    .io_tlbw_port_bits_entry_lo0_pfn(cp0_io_tlbw_port_bits_entry_lo0_pfn),
    .io_tlbw_port_bits_entry_lo0_c(cp0_io_tlbw_port_bits_entry_lo0_c),
    .io_tlbw_port_bits_entry_lo0_d(cp0_io_tlbw_port_bits_entry_lo0_d),
    .io_tlbw_port_bits_entry_lo0_v(cp0_io_tlbw_port_bits_entry_lo0_v),
    .io_tlbw_port_bits_entry_lo0_g(cp0_io_tlbw_port_bits_entry_lo0_g),
    .io_tlbw_port_bits_entry_lo1_pfn(cp0_io_tlbw_port_bits_entry_lo1_pfn),
    .io_tlbw_port_bits_entry_lo1_c(cp0_io_tlbw_port_bits_entry_lo1_c),
    .io_tlbw_port_bits_entry_lo1_d(cp0_io_tlbw_port_bits_entry_lo1_d),
    .io_tlbw_port_bits_entry_lo1_v(cp0_io_tlbw_port_bits_entry_lo1_v),
    .io_tlbw_port_bits_entry_lo1_g(cp0_io_tlbw_port_bits_entry_lo1_g),
    .io_tlbp_port_valid(cp0_io_tlbp_port_valid),
    .io_tlbp_port_bits_index_p(cp0_io_tlbp_port_bits_index_p),
    .io_tlbp_port_bits_index_index(cp0_io_tlbp_port_bits_index_index),
    .io_status_ERL(cp0_io_status_ERL),
    .io_ehu_valid(cp0_io_ehu_valid),
    .io_ehu_ip7(cp0_io_ehu_ip7),
    .io_ehu_ex_et(cp0_io_ehu_ex_et),
    .io_ehu_ex_code(cp0_io_ehu_ex_code),
    .io_ehu_ex_addr(cp0_io_ehu_ex_addr),
    .io_ehu_ex_asid(cp0_io_ehu_ex_asid),
    .io_ehu_wb_pc(cp0_io_ehu_wb_pc),
    .io_ehu_wb_is_ds(cp0_io_ehu_wb_is_ds),
    .io_ehu_wb_is_br(cp0_io_ehu_wb_is_br),
    .io_ehu_wb_npc(cp0_io_ehu_wb_npc),
    .io_ex_flush_valid(cp0_io_ex_flush_valid),
    .io_ex_flush_bits_br_target(cp0_io_ex_flush_bits_br_target)
  );
  TLB tlb ( // @[core.scala 30:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_iaddr_req_ready(tlb_io_iaddr_req_ready),
    .io_iaddr_req_valid(tlb_io_iaddr_req_valid),
    .io_iaddr_req_bits_vaddr(tlb_io_iaddr_req_bits_vaddr),
    .io_iaddr_resp_ready(tlb_io_iaddr_resp_ready),
    .io_iaddr_resp_valid(tlb_io_iaddr_resp_valid),
    .io_iaddr_resp_bits_paddr(tlb_io_iaddr_resp_bits_paddr),
    .io_iaddr_resp_bits_is_cached(tlb_io_iaddr_resp_bits_is_cached),
    .io_iaddr_resp_bits_ex_et(tlb_io_iaddr_resp_bits_ex_et),
    .io_iaddr_resp_bits_ex_code(tlb_io_iaddr_resp_bits_ex_code),
    .io_iaddr_resp_bits_ex_addr(tlb_io_iaddr_resp_bits_ex_addr),
    .io_iaddr_resp_bits_ex_asid(tlb_io_iaddr_resp_bits_ex_asid),
    .io_daddr_req_ready(tlb_io_daddr_req_ready),
    .io_daddr_req_valid(tlb_io_daddr_req_valid),
    .io_daddr_req_bits_func(tlb_io_daddr_req_bits_func),
    .io_daddr_req_bits_vaddr(tlb_io_daddr_req_bits_vaddr),
    .io_daddr_req_bits_len(tlb_io_daddr_req_bits_len),
    .io_daddr_req_bits_is_aligned(tlb_io_daddr_req_bits_is_aligned),
    .io_daddr_resp_bits_paddr(tlb_io_daddr_resp_bits_paddr),
    .io_daddr_resp_bits_ex_et(tlb_io_daddr_resp_bits_ex_et),
    .io_daddr_resp_bits_ex_code(tlb_io_daddr_resp_bits_ex_code),
    .io_daddr_resp_bits_ex_addr(tlb_io_daddr_resp_bits_ex_addr),
    .io_daddr_resp_bits_ex_asid(tlb_io_daddr_resp_bits_ex_asid),
    .io_rport_index(tlb_io_rport_index),
    .io_rport_entry_pagemask(tlb_io_rport_entry_pagemask),
    .io_rport_entry_vpn(tlb_io_rport_entry_vpn),
    .io_rport_entry_g(tlb_io_rport_entry_g),
    .io_rport_entry_asid(tlb_io_rport_entry_asid),
    .io_rport_entry_p0_pfn(tlb_io_rport_entry_p0_pfn),
    .io_rport_entry_p0_c(tlb_io_rport_entry_p0_c),
    .io_rport_entry_p0_d(tlb_io_rport_entry_p0_d),
    .io_rport_entry_p0_v(tlb_io_rport_entry_p0_v),
    .io_rport_entry_p1_pfn(tlb_io_rport_entry_p1_pfn),
    .io_rport_entry_p1_c(tlb_io_rport_entry_p1_c),
    .io_rport_entry_p1_d(tlb_io_rport_entry_p1_d),
    .io_rport_entry_p1_v(tlb_io_rport_entry_p1_v),
    .io_wport_valid(tlb_io_wport_valid),
    .io_wport_bits_index(tlb_io_wport_bits_index),
    .io_wport_bits_entry_pagemask(tlb_io_wport_bits_entry_pagemask),
    .io_wport_bits_entry_vpn(tlb_io_wport_bits_entry_vpn),
    .io_wport_bits_entry_g(tlb_io_wport_bits_entry_g),
    .io_wport_bits_entry_asid(tlb_io_wport_bits_entry_asid),
    .io_wport_bits_entry_p0_pfn(tlb_io_wport_bits_entry_p0_pfn),
    .io_wport_bits_entry_p0_c(tlb_io_wport_bits_entry_p0_c),
    .io_wport_bits_entry_p0_d(tlb_io_wport_bits_entry_p0_d),
    .io_wport_bits_entry_p0_v(tlb_io_wport_bits_entry_p0_v),
    .io_wport_bits_entry_p1_pfn(tlb_io_wport_bits_entry_p1_pfn),
    .io_wport_bits_entry_p1_c(tlb_io_wport_bits_entry_p1_c),
    .io_wport_bits_entry_p1_d(tlb_io_wport_bits_entry_p1_d),
    .io_wport_bits_entry_p1_v(tlb_io_wport_bits_entry_p1_v),
    .io_pport_entry_hi_vpn(tlb_io_pport_entry_hi_vpn),
    .io_pport_entry_hi_asid(tlb_io_pport_entry_hi_asid),
    .io_pport_index_p(tlb_io_pport_index_p),
    .io_pport_index_index(tlb_io_pport_index_index),
    .io_status_ERL(tlb_io_status_ERL),
    .io_br_flush_valid(tlb_io_br_flush_valid),
    .io_ex_flush_valid(tlb_io_ex_flush_valid)
  );
  MSU msu ( // @[core.scala 31:19]
    .clock(msu_clock),
    .reset(msu_reset),
    .io_fu_in_ready(msu_io_fu_in_ready),
    .io_fu_in_valid(msu_io_fu_in_valid),
    .io_fu_in_bits_wb_v(msu_io_fu_in_bits_wb_v),
    .io_fu_in_bits_wb_id(msu_io_fu_in_bits_wb_id),
    .io_fu_in_bits_wb_pc(msu_io_fu_in_bits_wb_pc),
    .io_fu_in_bits_wb_instr_op(msu_io_fu_in_bits_wb_instr_op),
    .io_fu_in_bits_wb_instr_rs_idx(msu_io_fu_in_bits_wb_instr_rs_idx),
    .io_fu_in_bits_wb_instr_rt_idx(msu_io_fu_in_bits_wb_instr_rt_idx),
    .io_fu_in_bits_wb_instr_rd_idx(msu_io_fu_in_bits_wb_instr_rd_idx),
    .io_fu_in_bits_wb_instr_shamt(msu_io_fu_in_bits_wb_instr_shamt),
    .io_fu_in_bits_wb_instr_func(msu_io_fu_in_bits_wb_instr_func),
    .io_fu_in_bits_wb_rd_idx(msu_io_fu_in_bits_wb_rd_idx),
    .io_fu_in_bits_wb_wen(msu_io_fu_in_bits_wb_wen),
    .io_fu_in_bits_wb_data(msu_io_fu_in_bits_wb_data),
    .io_fu_in_bits_wb_ip7(msu_io_fu_in_bits_wb_ip7),
    .io_fu_in_bits_wb_is_ds(msu_io_fu_in_bits_wb_is_ds),
    .io_fu_in_bits_wb_is_br(msu_io_fu_in_bits_wb_is_br),
    .io_fu_in_bits_wb_npc(msu_io_fu_in_bits_wb_npc),
    .io_fu_in_bits_ops_fu_type(msu_io_fu_in_bits_ops_fu_type),
    .io_fu_in_bits_ops_fu_op(msu_io_fu_in_bits_ops_fu_op),
    .io_fu_in_bits_ops_op1(msu_io_fu_in_bits_ops_op1),
    .io_fu_in_bits_ops_op2(msu_io_fu_in_bits_ops_op2),
    .io_fu_in_bits_is_cached(msu_io_fu_in_bits_is_cached),
    .io_wb_valid(msu_io_wb_valid),
    .io_wb_bits_v(msu_io_wb_bits_v),
    .io_wb_bits_id(msu_io_wb_bits_id),
    .io_wb_bits_pc(msu_io_wb_bits_pc),
    .io_wb_bits_instr_op(msu_io_wb_bits_instr_op),
    .io_wb_bits_instr_rs_idx(msu_io_wb_bits_instr_rs_idx),
    .io_wb_bits_instr_rt_idx(msu_io_wb_bits_instr_rt_idx),
    .io_wb_bits_instr_rd_idx(msu_io_wb_bits_instr_rd_idx),
    .io_wb_bits_instr_shamt(msu_io_wb_bits_instr_shamt),
    .io_wb_bits_instr_func(msu_io_wb_bits_instr_func),
    .io_wb_bits_rd_idx(msu_io_wb_bits_rd_idx),
    .io_wb_bits_wen(msu_io_wb_bits_wen),
    .io_wb_bits_data(msu_io_wb_bits_data),
    .io_wb_bits_ip7(msu_io_wb_bits_ip7),
    .io_divider_data_dividend_tvalid(msu_io_divider_data_dividend_tvalid),
    .io_divider_data_divisor_tvalid(msu_io_divider_data_divisor_tvalid),
    .io_divider_data_dout_tvalid(msu_io_divider_data_dout_tvalid),
    .io_divider_data_dividend_tdata(msu_io_divider_data_dividend_tdata),
    .io_divider_data_divisor_tdata(msu_io_divider_data_divisor_tdata),
    .io_divider_data_dout_tdata(msu_io_divider_data_dout_tdata),
    .io_multiplier_data_a(msu_io_multiplier_data_a),
    .io_multiplier_data_b(msu_io_multiplier_data_b),
    .io_multiplier_data_dout(msu_io_multiplier_data_dout),
    .io_dmem_req_ready(msu_io_dmem_req_ready),
    .io_dmem_req_valid(msu_io_dmem_req_valid),
    .io_dmem_req_bits_is_cached(msu_io_dmem_req_bits_is_cached),
    .io_dmem_req_bits_addr(msu_io_dmem_req_bits_addr),
    .io_dmem_req_bits_len(msu_io_dmem_req_bits_len),
    .io_dmem_req_bits_strb(msu_io_dmem_req_bits_strb),
    .io_dmem_req_bits_data(msu_io_dmem_req_bits_data),
    .io_dmem_req_bits_func(msu_io_dmem_req_bits_func),
    .io_dmem_resp_valid(msu_io_dmem_resp_valid),
    .io_dmem_resp_bits_data(msu_io_dmem_resp_bits_data)
  );
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[core.scala 73:15]
  assign io_imem_req_bits_is_cached = ifu_io_imem_req_bits_is_cached; // @[core.scala 73:15]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[core.scala 73:15]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[core.scala 73:15]
  assign io_dmem_req_valid = msu_io_dmem_req_valid; // @[core.scala 74:15]
  assign io_dmem_req_bits_is_cached = msu_io_dmem_req_bits_is_cached; // @[core.scala 74:15]
  assign io_dmem_req_bits_addr = msu_io_dmem_req_bits_addr; // @[core.scala 74:15]
  assign io_dmem_req_bits_len = msu_io_dmem_req_bits_len; // @[core.scala 74:15]
  assign io_dmem_req_bits_strb = msu_io_dmem_req_bits_strb; // @[core.scala 74:15]
  assign io_dmem_req_bits_data = msu_io_dmem_req_bits_data; // @[core.scala 74:15]
  assign io_dmem_req_bits_func = msu_io_dmem_req_bits_func; // @[core.scala 74:15]
  assign io_icache_control_valid = exu_io_icache_control_valid; // @[core.scala 96:21]
  assign io_icache_control_bits_op = exu_io_icache_control_bits_op; // @[core.scala 96:21]
  assign io_icache_control_bits_addr = exu_io_icache_control_bits_addr; // @[core.scala 96:21]
  assign io_commit_valid = rf_io_commit_valid; // @[core.scala 77:13]
  assign io_commit_pc = rf_io_commit_pc; // @[core.scala 77:13]
  assign io_commit_instr = rf_io_commit_instr; // @[core.scala 77:13]
  assign io_commit_ip7 = rf_io_commit_ip7; // @[core.scala 77:13]
  assign io_commit_gpr_0 = rf_io_commit_gpr_0; // @[core.scala 77:13]
  assign io_commit_gpr_1 = rf_io_commit_gpr_1; // @[core.scala 77:13]
  assign io_commit_gpr_2 = rf_io_commit_gpr_2; // @[core.scala 77:13]
  assign io_commit_gpr_3 = rf_io_commit_gpr_3; // @[core.scala 77:13]
  assign io_commit_gpr_4 = rf_io_commit_gpr_4; // @[core.scala 77:13]
  assign io_commit_gpr_5 = rf_io_commit_gpr_5; // @[core.scala 77:13]
  assign io_commit_gpr_6 = rf_io_commit_gpr_6; // @[core.scala 77:13]
  assign io_commit_gpr_7 = rf_io_commit_gpr_7; // @[core.scala 77:13]
  assign io_commit_gpr_8 = rf_io_commit_gpr_8; // @[core.scala 77:13]
  assign io_commit_gpr_9 = rf_io_commit_gpr_9; // @[core.scala 77:13]
  assign io_commit_gpr_10 = rf_io_commit_gpr_10; // @[core.scala 77:13]
  assign io_commit_gpr_11 = rf_io_commit_gpr_11; // @[core.scala 77:13]
  assign io_commit_gpr_12 = rf_io_commit_gpr_12; // @[core.scala 77:13]
  assign io_commit_gpr_13 = rf_io_commit_gpr_13; // @[core.scala 77:13]
  assign io_commit_gpr_14 = rf_io_commit_gpr_14; // @[core.scala 77:13]
  assign io_commit_gpr_15 = rf_io_commit_gpr_15; // @[core.scala 77:13]
  assign io_commit_gpr_16 = rf_io_commit_gpr_16; // @[core.scala 77:13]
  assign io_commit_gpr_17 = rf_io_commit_gpr_17; // @[core.scala 77:13]
  assign io_commit_gpr_18 = rf_io_commit_gpr_18; // @[core.scala 77:13]
  assign io_commit_gpr_19 = rf_io_commit_gpr_19; // @[core.scala 77:13]
  assign io_commit_gpr_20 = rf_io_commit_gpr_20; // @[core.scala 77:13]
  assign io_commit_gpr_21 = rf_io_commit_gpr_21; // @[core.scala 77:13]
  assign io_commit_gpr_22 = rf_io_commit_gpr_22; // @[core.scala 77:13]
  assign io_commit_gpr_23 = rf_io_commit_gpr_23; // @[core.scala 77:13]
  assign io_commit_gpr_24 = rf_io_commit_gpr_24; // @[core.scala 77:13]
  assign io_commit_gpr_25 = rf_io_commit_gpr_25; // @[core.scala 77:13]
  assign io_commit_gpr_26 = rf_io_commit_gpr_26; // @[core.scala 77:13]
  assign io_commit_gpr_27 = rf_io_commit_gpr_27; // @[core.scala 77:13]
  assign io_commit_gpr_28 = rf_io_commit_gpr_28; // @[core.scala 77:13]
  assign io_commit_gpr_29 = rf_io_commit_gpr_29; // @[core.scala 77:13]
  assign io_commit_gpr_30 = rf_io_commit_gpr_30; // @[core.scala 77:13]
  assign io_commit_gpr_31 = rf_io_commit_gpr_31; // @[core.scala 77:13]
  assign io_commit_rd_idx = rf_io_commit_rd_idx; // @[core.scala 77:13]
  assign io_commit_wdata = rf_io_commit_wdata; // @[core.scala 77:13]
  assign io_commit_wen = rf_io_commit_wen; // @[core.scala 77:13]
  assign io_br_flush = idu_io_br_flush_valid; // @[core.scala 80:15]
  assign io_ex_flush = cp0_io_ex_flush_valid; // @[core.scala 81:15]
  assign io_multiplier_data_a = msu_io_multiplier_data_a; // @[core.scala 93:21]
  assign io_multiplier_data_b = msu_io_multiplier_data_b; // @[core.scala 93:21]
  assign io_divider_data_dividend_tvalid = msu_io_divider_data_dividend_tvalid; // @[core.scala 94:18]
  assign io_divider_data_divisor_tvalid = msu_io_divider_data_divisor_tvalid; // @[core.scala 94:18]
  assign io_divider_data_dividend_tdata = msu_io_divider_data_dividend_tdata; // @[core.scala 94:18]
  assign io_divider_data_divisor_tdata = msu_io_divider_data_divisor_tdata; // @[core.scala 94:18]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_bp_valid = exu_io_bp_valid; // @[core.scala 55:13]
  assign rf_io_bp_bits_v = exu_io_bp_bits_v; // @[core.scala 55:13]
  assign rf_io_bp_bits_rd_idx = exu_io_bp_bits_rd_idx; // @[core.scala 55:13]
  assign rf_io_bp_bits_wen = exu_io_bp_bits_wen; // @[core.scala 55:13]
  assign rf_io_bp_bits_data = exu_io_bp_bits_data; // @[core.scala 55:13]
  assign rf_io_wb_valid = msu_io_wb_valid; // @[core.scala 53:13]
  assign rf_io_wb_bits_v = msu_io_wb_bits_v; // @[core.scala 53:13]
  assign rf_io_wb_bits_id = msu_io_wb_bits_id; // @[core.scala 53:13]
  assign rf_io_wb_bits_pc = msu_io_wb_bits_pc; // @[core.scala 53:13]
  assign rf_io_wb_bits_instr_op = msu_io_wb_bits_instr_op; // @[core.scala 53:13]
  assign rf_io_wb_bits_instr_rs_idx = msu_io_wb_bits_instr_rs_idx; // @[core.scala 53:13]
  assign rf_io_wb_bits_instr_rt_idx = msu_io_wb_bits_instr_rt_idx; // @[core.scala 53:13]
  assign rf_io_wb_bits_instr_rd_idx = msu_io_wb_bits_instr_rd_idx; // @[core.scala 53:13]
  assign rf_io_wb_bits_instr_shamt = msu_io_wb_bits_instr_shamt; // @[core.scala 53:13]
  assign rf_io_wb_bits_instr_func = msu_io_wb_bits_instr_func; // @[core.scala 53:13]
  assign rf_io_wb_bits_rd_idx = msu_io_wb_bits_rd_idx; // @[core.scala 53:13]
  assign rf_io_wb_bits_wen = msu_io_wb_bits_wen; // @[core.scala 53:13]
  assign rf_io_wb_bits_data = msu_io_wb_bits_data; // @[core.scala 53:13]
  assign rf_io_wb_bits_ip7 = msu_io_wb_bits_ip7; // @[core.scala 53:13]
  assign rf_io_rfio_rs_idx = idu_io_rfio_rs_idx; // @[core.scala 56:15]
  assign rf_io_rfio_rt_idx = idu_io_rfio_rt_idx; // @[core.scala 56:15]
  assign rf_io_rfio_wen = idu_io_rfio_wen; // @[core.scala 56:15]
  assign rf_io_rfio_wid = idu_io_rfio_wid; // @[core.scala 56:15]
  assign rf_io_rfio_rd_idx = idu_io_rfio_rd_idx; // @[core.scala 56:15]
  assign rf_io_ex_flush_valid = cp0_io_ex_flush_valid; // @[core.scala 87:18]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[core.scala 73:15]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[core.scala 73:15]
  assign ifu_io_imem_resp_bits_data = io_imem_resp_bits_data; // @[core.scala 73:15]
  assign ifu_io_iaddr_req_ready = tlb_io_iaddr_req_ready; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_valid = tlb_io_iaddr_resp_valid; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_bits_paddr = tlb_io_iaddr_resp_bits_paddr; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_bits_is_cached = tlb_io_iaddr_resp_bits_is_cached; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_bits_ex_et = tlb_io_iaddr_resp_bits_ex_et; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_bits_ex_code = tlb_io_iaddr_resp_bits_ex_code; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_bits_ex_addr = tlb_io_iaddr_resp_bits_ex_addr; // @[core.scala 63:16]
  assign ifu_io_iaddr_resp_bits_ex_asid = tlb_io_iaddr_resp_bits_ex_asid; // @[core.scala 63:16]
  assign ifu_io_fu_out_ready = idu_io_fu_in_ready; // @[core.scala 44:17]
  assign ifu_io_br_flush_valid = idu_io_br_flush_valid; // @[core.scala 82:19]
  assign ifu_io_br_flush_bits_br_target = idu_io_br_flush_bits_br_target; // @[core.scala 82:19]
  assign ifu_io_ex_flush_valid = cp0_io_ex_flush_valid; // @[core.scala 83:19]
  assign ifu_io_ex_flush_bits_br_target = cp0_io_ex_flush_bits_br_target; // @[core.scala 83:19]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_fu_in_valid = ifu_io_fu_out_valid; // @[core.scala 44:17]
  assign idu_io_fu_in_bits_pc = ifu_io_fu_out_bits_pc; // @[core.scala 44:17]
  assign idu_io_fu_in_bits_instr = ifu_io_fu_out_bits_instr; // @[core.scala 44:17]
  assign idu_io_fu_in_bits_ex_et = ifu_io_fu_out_bits_ex_et; // @[core.scala 44:17]
  assign idu_io_fu_in_bits_ex_code = ifu_io_fu_out_bits_ex_code; // @[core.scala 44:17]
  assign idu_io_fu_in_bits_ex_addr = ifu_io_fu_out_bits_ex_addr; // @[core.scala 44:17]
  assign idu_io_fu_in_bits_ex_asid = ifu_io_fu_out_bits_ex_asid; // @[core.scala 44:17]
  assign idu_io_fu_out_ready = exu_io_fu_in_ready; // @[core.scala 45:17]
  assign idu_io_rfio_rs_data_valid = rf_io_rfio_rs_data_valid; // @[core.scala 56:15]
  assign idu_io_rfio_rs_data_bits = rf_io_rfio_rs_data_bits; // @[core.scala 56:15]
  assign idu_io_rfio_rt_data_valid = rf_io_rfio_rt_data_valid; // @[core.scala 56:15]
  assign idu_io_rfio_rt_data_bits = rf_io_rfio_rt_data_bits; // @[core.scala 56:15]
  assign idu_io_ex_flush_valid = cp0_io_ex_flush_valid; // @[core.scala 84:19]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_fu_in_valid = idu_io_fu_out_valid; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_v = idu_io_fu_out_bits_wb_v; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_id = idu_io_fu_out_bits_wb_id; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_pc = idu_io_fu_out_bits_wb_pc; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_instr_op = idu_io_fu_out_bits_wb_instr_op; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_instr_rs_idx = idu_io_fu_out_bits_wb_instr_rs_idx; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_instr_rt_idx = idu_io_fu_out_bits_wb_instr_rt_idx; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_instr_rd_idx = idu_io_fu_out_bits_wb_instr_rd_idx; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_instr_shamt = idu_io_fu_out_bits_wb_instr_shamt; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_instr_func = idu_io_fu_out_bits_wb_instr_func; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_rd_idx = idu_io_fu_out_bits_wb_rd_idx; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_wen = idu_io_fu_out_bits_wb_wen; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_data = idu_io_fu_out_bits_wb_data; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_is_ds = idu_io_fu_out_bits_wb_is_ds; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_is_br = idu_io_fu_out_bits_wb_is_br; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_wb_npc = idu_io_fu_out_bits_wb_npc; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ops_fu_type = idu_io_fu_out_bits_ops_fu_type; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ops_fu_op = idu_io_fu_out_bits_ops_fu_op; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ops_op1 = idu_io_fu_out_bits_ops_op1; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ops_op2 = idu_io_fu_out_bits_ops_op2; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ex_et = idu_io_fu_out_bits_ex_et; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ex_code = idu_io_fu_out_bits_ex_code; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ex_addr = idu_io_fu_out_bits_ex_addr; // @[core.scala 45:17]
  assign exu_io_fu_in_bits_ex_asid = idu_io_fu_out_bits_ex_asid; // @[core.scala 45:17]
  assign exu_io_fu_out_ready = ehu_io_fu_in_ready; // @[core.scala 46:17]
  assign exu_io_cp0_rport_data = cp0_io_rport_data; // @[core.scala 59:20]
  assign exu_io_cp0_tlbr_port_index_index = cp0_io_tlbr_port_index_index; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_pagemask_mask = cp0_io_tlbr_port_pagemask_mask; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_hi_vpn = cp0_io_tlbr_port_entry_hi_vpn; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_hi_asid = cp0_io_tlbr_port_entry_hi_asid; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo0_pfn = cp0_io_tlbr_port_entry_lo0_pfn; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo0_c = cp0_io_tlbr_port_entry_lo0_c; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo0_d = cp0_io_tlbr_port_entry_lo0_d; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo0_v = cp0_io_tlbr_port_entry_lo0_v; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo0_g = cp0_io_tlbr_port_entry_lo0_g; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo1_pfn = cp0_io_tlbr_port_entry_lo1_pfn; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo1_c = cp0_io_tlbr_port_entry_lo1_c; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo1_d = cp0_io_tlbr_port_entry_lo1_d; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo1_v = cp0_io_tlbr_port_entry_lo1_v; // @[core.scala 65:24]
  assign exu_io_cp0_tlbr_port_entry_lo1_g = cp0_io_tlbr_port_entry_lo1_g; // @[core.scala 65:24]
  assign exu_io_daddr_resp_bits_paddr = tlb_io_daddr_resp_bits_paddr; // @[core.scala 64:16]
  assign exu_io_daddr_resp_bits_ex_et = tlb_io_daddr_resp_bits_ex_et; // @[core.scala 64:16]
  assign exu_io_daddr_resp_bits_ex_code = tlb_io_daddr_resp_bits_ex_code; // @[core.scala 64:16]
  assign exu_io_daddr_resp_bits_ex_addr = tlb_io_daddr_resp_bits_ex_addr; // @[core.scala 64:16]
  assign exu_io_daddr_resp_bits_ex_asid = tlb_io_daddr_resp_bits_ex_asid; // @[core.scala 64:16]
  assign exu_io_tlb_rport_entry_pagemask = tlb_io_rport_entry_pagemask; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_vpn = tlb_io_rport_entry_vpn; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_g = tlb_io_rport_entry_g; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_asid = tlb_io_rport_entry_asid; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p0_pfn = tlb_io_rport_entry_p0_pfn; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p0_c = tlb_io_rport_entry_p0_c; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p0_d = tlb_io_rport_entry_p0_d; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p0_v = tlb_io_rport_entry_p0_v; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p1_pfn = tlb_io_rport_entry_p1_pfn; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p1_c = tlb_io_rport_entry_p1_c; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p1_d = tlb_io_rport_entry_p1_d; // @[core.scala 68:20]
  assign exu_io_tlb_rport_entry_p1_v = tlb_io_rport_entry_p1_v; // @[core.scala 68:20]
  assign exu_io_tlb_pport_index_p = tlb_io_pport_index_p; // @[core.scala 70:20]
  assign exu_io_tlb_pport_index_index = tlb_io_pport_index_index; // @[core.scala 70:20]
  assign exu_io_ex_flush_valid = cp0_io_ex_flush_valid; // @[core.scala 85:19]
  assign ehu_clock = clock;
  assign ehu_reset = reset;
  assign ehu_io_fu_in_valid = exu_io_fu_out_valid; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_v = exu_io_fu_out_bits_wb_v; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_id = exu_io_fu_out_bits_wb_id; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_pc = exu_io_fu_out_bits_wb_pc; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_instr_op = exu_io_fu_out_bits_wb_instr_op; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_instr_rs_idx = exu_io_fu_out_bits_wb_instr_rs_idx; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_instr_rt_idx = exu_io_fu_out_bits_wb_instr_rt_idx; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_instr_rd_idx = exu_io_fu_out_bits_wb_instr_rd_idx; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_instr_shamt = exu_io_fu_out_bits_wb_instr_shamt; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_instr_func = exu_io_fu_out_bits_wb_instr_func; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_rd_idx = exu_io_fu_out_bits_wb_rd_idx; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_wen = exu_io_fu_out_bits_wb_wen; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_data = exu_io_fu_out_bits_wb_data; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_is_ds = exu_io_fu_out_bits_wb_is_ds; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_is_br = exu_io_fu_out_bits_wb_is_br; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_wb_npc = exu_io_fu_out_bits_wb_npc; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ops_fu_type = exu_io_fu_out_bits_ops_fu_type; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ops_fu_op = exu_io_fu_out_bits_ops_fu_op; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ops_op1 = exu_io_fu_out_bits_ops_op1; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ops_op2 = exu_io_fu_out_bits_ops_op2; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ex_et = exu_io_fu_out_bits_ex_et; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ex_code = exu_io_fu_out_bits_ex_code; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ex_addr = exu_io_fu_out_bits_ex_addr; // @[core.scala 46:17]
  assign ehu_io_fu_in_bits_ex_asid = exu_io_fu_out_bits_ex_asid; // @[core.scala 46:17]
  assign ehu_io_fu_out_ready = msu_io_fu_in_ready; // @[core.scala 47:17]
  assign ehu_io_cp0_ip7 = cp0_io_ehu_ip7; // @[core.scala 50:14]
  assign ehu_io_ex_flush_valid = cp0_io_ex_flush_valid; // @[core.scala 86:19]
  assign cp0_clock = clock;
  assign cp0_reset = reset;
  assign cp0_io_rport_addr = exu_io_cp0_rport_addr; // @[core.scala 59:20]
  assign cp0_io_wport_valid = exu_io_cp0_wport_valid; // @[core.scala 60:20]
  assign cp0_io_wport_bits_addr = exu_io_cp0_wport_bits_addr; // @[core.scala 60:20]
  assign cp0_io_wport_bits_data = exu_io_cp0_wport_bits_data; // @[core.scala 60:20]
  assign cp0_io_tlbw_port_valid = exu_io_cp0_tlbw_port_valid; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_pagemask_mask = exu_io_cp0_tlbw_port_bits_pagemask_mask; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_hi_vpn = exu_io_cp0_tlbw_port_bits_entry_hi_vpn; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_hi_asid = exu_io_cp0_tlbw_port_bits_entry_hi_asid; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo0_pfn = exu_io_cp0_tlbw_port_bits_entry_lo0_pfn; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo0_c = exu_io_cp0_tlbw_port_bits_entry_lo0_c; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo0_d = exu_io_cp0_tlbw_port_bits_entry_lo0_d; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo0_v = exu_io_cp0_tlbw_port_bits_entry_lo0_v; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo0_g = exu_io_cp0_tlbw_port_bits_entry_lo0_g; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo1_pfn = exu_io_cp0_tlbw_port_bits_entry_lo1_pfn; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo1_c = exu_io_cp0_tlbw_port_bits_entry_lo1_c; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo1_d = exu_io_cp0_tlbw_port_bits_entry_lo1_d; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo1_v = exu_io_cp0_tlbw_port_bits_entry_lo1_v; // @[core.scala 66:24]
  assign cp0_io_tlbw_port_bits_entry_lo1_g = exu_io_cp0_tlbw_port_bits_entry_lo1_g; // @[core.scala 66:24]
  assign cp0_io_tlbp_port_valid = exu_io_cp0_tlbp_port_valid; // @[core.scala 67:24]
  assign cp0_io_tlbp_port_bits_index_p = exu_io_cp0_tlbp_port_bits_index_p; // @[core.scala 67:24]
  assign cp0_io_tlbp_port_bits_index_index = exu_io_cp0_tlbp_port_bits_index_index; // @[core.scala 67:24]
  assign cp0_io_ehu_valid = ehu_io_cp0_valid; // @[core.scala 50:14]
  assign cp0_io_ehu_ex_et = ehu_io_cp0_ex_et; // @[core.scala 50:14]
  assign cp0_io_ehu_ex_code = ehu_io_cp0_ex_code; // @[core.scala 50:14]
  assign cp0_io_ehu_ex_addr = ehu_io_cp0_ex_addr; // @[core.scala 50:14]
  assign cp0_io_ehu_ex_asid = ehu_io_cp0_ex_asid; // @[core.scala 50:14]
  assign cp0_io_ehu_wb_pc = ehu_io_cp0_wb_pc; // @[core.scala 50:14]
  assign cp0_io_ehu_wb_is_ds = ehu_io_cp0_wb_is_ds; // @[core.scala 50:14]
  assign cp0_io_ehu_wb_is_br = ehu_io_cp0_wb_is_br; // @[core.scala 50:14]
  assign cp0_io_ehu_wb_npc = ehu_io_cp0_wb_npc; // @[core.scala 50:14]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_iaddr_req_valid = ifu_io_iaddr_req_valid; // @[core.scala 63:16]
  assign tlb_io_iaddr_req_bits_vaddr = ifu_io_iaddr_req_bits_vaddr; // @[core.scala 63:16]
  assign tlb_io_iaddr_resp_ready = ifu_io_iaddr_resp_ready; // @[core.scala 63:16]
  assign tlb_io_daddr_req_valid = exu_io_daddr_req_valid; // @[core.scala 64:16]
  assign tlb_io_daddr_req_bits_func = exu_io_daddr_req_bits_func; // @[core.scala 64:16]
  assign tlb_io_daddr_req_bits_vaddr = exu_io_daddr_req_bits_vaddr; // @[core.scala 64:16]
  assign tlb_io_daddr_req_bits_len = exu_io_daddr_req_bits_len; // @[core.scala 64:16]
  assign tlb_io_daddr_req_bits_is_aligned = exu_io_daddr_req_bits_is_aligned; // @[core.scala 64:16]
  assign tlb_io_rport_index = exu_io_tlb_rport_index; // @[core.scala 68:20]
  assign tlb_io_wport_valid = exu_io_tlb_wport_valid; // @[core.scala 69:20]
  assign tlb_io_wport_bits_index = exu_io_tlb_wport_bits_index; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_pagemask = exu_io_tlb_wport_bits_entry_pagemask; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_vpn = exu_io_tlb_wport_bits_entry_vpn; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_g = exu_io_tlb_wport_bits_entry_g; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_asid = exu_io_tlb_wport_bits_entry_asid; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p0_pfn = exu_io_tlb_wport_bits_entry_p0_pfn; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p0_c = exu_io_tlb_wport_bits_entry_p0_c; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p0_d = exu_io_tlb_wport_bits_entry_p0_d; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p0_v = exu_io_tlb_wport_bits_entry_p0_v; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p1_pfn = exu_io_tlb_wport_bits_entry_p1_pfn; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p1_c = exu_io_tlb_wport_bits_entry_p1_c; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p1_d = exu_io_tlb_wport_bits_entry_p1_d; // @[core.scala 69:20]
  assign tlb_io_wport_bits_entry_p1_v = exu_io_tlb_wport_bits_entry_p1_v; // @[core.scala 69:20]
  assign tlb_io_pport_entry_hi_vpn = exu_io_tlb_pport_entry_hi_vpn; // @[core.scala 70:20]
  assign tlb_io_pport_entry_hi_asid = exu_io_tlb_pport_entry_hi_asid; // @[core.scala 70:20]
  assign tlb_io_status_ERL = cp0_io_status_ERL; // @[core.scala 91:17]
  assign tlb_io_br_flush_valid = idu_io_br_flush_valid; // @[core.scala 88:19]
  assign tlb_io_ex_flush_valid = cp0_io_ex_flush_valid; // @[core.scala 89:19]
  assign msu_clock = clock;
  assign msu_reset = reset;
  assign msu_io_fu_in_valid = ehu_io_fu_out_valid; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_v = ehu_io_fu_out_bits_wb_v; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_id = ehu_io_fu_out_bits_wb_id; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_pc = ehu_io_fu_out_bits_wb_pc; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_instr_op = ehu_io_fu_out_bits_wb_instr_op; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_instr_rs_idx = ehu_io_fu_out_bits_wb_instr_rs_idx; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_instr_rt_idx = ehu_io_fu_out_bits_wb_instr_rt_idx; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_instr_rd_idx = ehu_io_fu_out_bits_wb_instr_rd_idx; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_instr_shamt = ehu_io_fu_out_bits_wb_instr_shamt; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_instr_func = ehu_io_fu_out_bits_wb_instr_func; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_rd_idx = ehu_io_fu_out_bits_wb_rd_idx; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_wen = ehu_io_fu_out_bits_wb_wen; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_data = ehu_io_fu_out_bits_wb_data; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_ip7 = ehu_io_fu_out_bits_wb_ip7; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_is_ds = ehu_io_fu_out_bits_wb_is_ds; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_is_br = ehu_io_fu_out_bits_wb_is_br; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_wb_npc = ehu_io_fu_out_bits_wb_npc; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_ops_fu_type = ehu_io_fu_out_bits_ops_fu_type; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_ops_fu_op = ehu_io_fu_out_bits_ops_fu_op; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_ops_op1 = ehu_io_fu_out_bits_ops_op1; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_ops_op2 = ehu_io_fu_out_bits_ops_op2; // @[core.scala 47:17]
  assign msu_io_fu_in_bits_is_cached = ehu_io_fu_out_bits_is_cached; // @[core.scala 47:17]
  assign msu_io_divider_data_dout_tvalid = io_divider_data_dout_tvalid; // @[core.scala 94:18]
  assign msu_io_divider_data_dout_tdata = io_divider_data_dout_tdata; // @[core.scala 94:18]
  assign msu_io_multiplier_data_dout = io_multiplier_data_dout; // @[core.scala 93:21]
  assign msu_io_dmem_req_ready = io_dmem_req_ready; // @[core.scala 74:15]
  assign msu_io_dmem_resp_valid = io_dmem_resp_valid; // @[core.scala 74:15]
  assign msu_io_dmem_resp_bits_data = io_dmem_resp_bits_data; // @[core.scala 74:15]
endmodule
module CrossbarNx1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input         io_in_0_req_bits_is_cached,
  input  [31:0] io_in_0_req_bits_addr,
  input  [1:0]  io_in_0_req_bits_len,
  input  [3:0]  io_in_0_req_bits_strb,
  output        io_in_0_resp_valid,
  output [31:0] io_in_0_resp_bits_data,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input         io_in_1_req_bits_is_cached,
  input  [31:0] io_in_1_req_bits_addr,
  input  [1:0]  io_in_1_req_bits_len,
  input  [3:0]  io_in_1_req_bits_strb,
  input  [31:0] io_in_1_req_bits_data,
  input         io_in_1_req_bits_func,
  output        io_in_1_resp_valid,
  output [31:0] io_in_1_resp_bits_data,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output        io_out_req_bits_is_cached,
  output [31:0] io_out_req_bits_addr,
  output [1:0]  io_out_req_bits_len,
  output [3:0]  io_out_req_bits_strb,
  output [31:0] io_out_req_bits_data,
  output        io_out_req_bits_func,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [31:0] io_out_resp_bits_data
);
  reg [1:0] q_datas [0:2]; // @[bridge.scala 145:20]
  reg [31:0] _RAND_0;
  wire [1:0] q_datas_q_out_data; // @[bridge.scala 145:20]
  wire [1:0] q_datas_q_out_addr; // @[bridge.scala 145:20]
  reg [31:0] _RAND_1;
  wire [1:0] q_datas__T_61_data; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_61_addr; // @[bridge.scala 145:20]
  reg [31:0] _RAND_2;
  wire [1:0] q_datas__T_63_data; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_63_addr; // @[bridge.scala 145:20]
  reg [31:0] _RAND_3;
  wire [1:0] q_datas__T_60_data; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_60_addr; // @[bridge.scala 145:20]
  wire  q_datas__T_60_mask; // @[bridge.scala 145:20]
  wire  q_datas__T_60_en; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_62_data; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_62_addr; // @[bridge.scala 145:20]
  wire  q_datas__T_62_mask; // @[bridge.scala 145:20]
  wire  q_datas__T_62_en; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_64_data; // @[bridge.scala 145:20]
  wire [1:0] q_datas__T_64_addr; // @[bridge.scala 145:20]
  wire  q_datas__T_64_mask; // @[bridge.scala 145:20]
  wire  q_datas__T_64_en; // @[bridge.scala 145:20]
  wire [1:0] _T = {io_in_0_req_valid,io_in_1_req_valid}; // @[Cat.scala 29:58]
  wire [1:0] in_valids = {_T[0],_T[1]}; // @[Cat.scala 29:58]
  reg [30:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  wire  _T_10 = value == 31'h7ffffffe; // @[Counter.scala 38:24]
  wire [30:0] _T_12 = value + 31'h1; // @[Counter.scala 39:22]
  wire  _T_17 = ~in_valids[0]; // @[utils.scala 111:21]
  wire  _T_18 = in_valids[1] & _T_17; // @[utils.scala 111:18]
  wire [1:0] _T_20 = {_T_18,in_valids[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_23 = {in_valids[0],in_valids[1]}; // @[Cat.scala 29:58]
  wire  _T_27 = ~_T_23[0]; // @[utils.scala 111:21]
  wire  _T_28 = _T_23[1] & _T_27; // @[utils.scala 111:18]
  wire [1:0] _T_30 = {_T_28,_T_23[0]}; // @[Cat.scala 29:58]
  wire [1:0] _T_33 = {_T_30[0],_T_30[1]}; // @[Cat.scala 29:58]
  wire [1:0] in_valids_1H = value[0] ? _T_20 : _T_33; // @[bridge.scala 138:25]
  wire [71:0] _T_40 = {io_in_0_req_bits_is_cached,io_in_0_req_bits_addr,io_in_0_req_bits_len,io_in_0_req_bits_strb,32'h0,1'h0}; // @[Mux.scala 27:72]
  wire [71:0] _T_41 = in_valids_1H[0] ? _T_40 : 72'h0; // @[Mux.scala 27:72]
  wire [71:0] _T_46 = {io_in_1_req_bits_is_cached,io_in_1_req_bits_addr,io_in_1_req_bits_len,io_in_1_req_bits_strb,io_in_1_req_bits_data,io_in_1_req_bits_func}; // @[Mux.scala 27:72]
  wire [71:0] _T_47 = in_valids_1H[1] ? _T_46 : 72'h0; // @[Mux.scala 27:72]
  wire [71:0] _T_48 = _T_41 | _T_47; // @[Mux.scala 27:72]
  reg [1:0] q_data_sz; // @[bridge.scala 144:26]
  reg [31:0] _RAND_5;
  wire  _T_59 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_11 = {{1'd0}, _T_59}; // @[bridge.scala 153:26]
  wire [1:0] _T_67 = q_data_sz + _GEN_11; // @[bridge.scala 153:26]
  wire  _T_68 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _GEN_12 = {{1'd0}, _T_68}; // @[bridge.scala 153:46]
  wire [1:0] _T_70 = _T_67 - _GEN_12; // @[bridge.scala 153:46]
  wire [1:0] _T_79 = q_datas_q_out_data; // @[bridge.scala 161:31]
  wire [1:0] _T_82 = ~q_data_sz; // @[bridge.scala 168:12]
  wire  _T_83 = _T_82 != 2'h0; // @[bridge.scala 168:24]
  wire  _T_85 = ~io_out_resp_valid; // @[bridge.scala 168:39]
  wire  _T_86 = _T_83 | _T_85; // @[bridge.scala 168:36]
  wire  _T_88 = _T_86 | reset; // @[bridge.scala 168:10]
  wire  _T_89 = ~_T_88; // @[bridge.scala 168:10]
  assign q_datas_q_out_addr = q_data_sz;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign q_datas_q_out_data = q_datas[q_datas_q_out_addr]; // @[bridge.scala 145:20]
  `else
  assign q_datas_q_out_data = q_datas_q_out_addr >= 2'h3 ? _RAND_1[1:0] : q_datas[q_datas_q_out_addr]; // @[bridge.scala 145:20]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign q_datas__T_61_addr = 2'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign q_datas__T_61_data = q_datas[q_datas__T_61_addr]; // @[bridge.scala 145:20]
  `else
  assign q_datas__T_61_data = q_datas__T_61_addr >= 2'h3 ? _RAND_2[1:0] : q_datas[q_datas__T_61_addr]; // @[bridge.scala 145:20]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign q_datas__T_63_addr = 2'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign q_datas__T_63_data = q_datas[q_datas__T_63_addr]; // @[bridge.scala 145:20]
  `else
  assign q_datas__T_63_data = q_datas__T_63_addr >= 2'h3 ? _RAND_3[1:0] : q_datas[q_datas__T_63_addr]; // @[bridge.scala 145:20]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign q_datas__T_60_data = q_datas__T_61_data;
  assign q_datas__T_60_addr = 2'h1;
  assign q_datas__T_60_mask = 1'h1;
  assign q_datas__T_60_en = io_out_req_ready & io_out_req_valid;
  assign q_datas__T_62_data = q_datas__T_63_data;
  assign q_datas__T_62_addr = 2'h2;
  assign q_datas__T_62_mask = 1'h1;
  assign q_datas__T_62_en = io_out_req_ready & io_out_req_valid;
  assign q_datas__T_64_data = value[0] ? _T_20 : _T_33;
  assign q_datas__T_64_addr = 2'h0;
  assign q_datas__T_64_mask = 1'h1;
  assign q_datas__T_64_en = io_out_req_ready & io_out_req_valid;
  assign io_in_0_req_ready = io_out_req_ready & in_valids_1H[0]; // @[bridge.scala 156:24]
  assign io_in_0_resp_valid = io_out_resp_valid & q_datas_q_out_data[0]; // @[bridge.scala 157:25]
  assign io_in_0_resp_bits_data = io_out_resp_bits_data; // @[bridge.scala 158:24]
  assign io_in_1_req_ready = io_out_req_ready & in_valids_1H[1]; // @[bridge.scala 156:24]
  assign io_in_1_resp_valid = io_out_resp_valid & q_datas_q_out_data[1]; // @[bridge.scala 157:25]
  assign io_in_1_resp_bits_data = io_out_resp_bits_data; // @[bridge.scala 158:24]
  assign io_out_req_valid = in_valids != 2'h0; // @[bridge.scala 162:20]
  assign io_out_req_bits_is_cached = _T_48[71]; // @[bridge.scala 163:19]
  assign io_out_req_bits_addr = _T_48[70:39]; // @[bridge.scala 163:19]
  assign io_out_req_bits_len = _T_48[38:37]; // @[bridge.scala 163:19]
  assign io_out_req_bits_strb = _T_48[36:33]; // @[bridge.scala 163:19]
  assign io_out_req_bits_data = _T_48[32:1]; // @[bridge.scala 163:19]
  assign io_out_req_bits_func = _T_48[0]; // @[bridge.scala 163:19]
  assign io_out_resp_ready = _T_79 != 2'h0; // @[bridge.scala 161:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    q_datas[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  _RAND_2 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  q_data_sz = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(q_datas__T_60_en & q_datas__T_60_mask) begin
      q_datas[q_datas__T_60_addr] <= q_datas__T_60_data; // @[bridge.scala 145:20]
    end
    if(q_datas__T_62_en & q_datas__T_62_mask) begin
      q_datas[q_datas__T_62_addr] <= q_datas__T_62_data; // @[bridge.scala 145:20]
    end
    if(q_datas__T_64_en & q_datas__T_64_mask) begin
      q_datas[q_datas__T_64_addr] <= q_datas__T_64_data; // @[bridge.scala 145:20]
    end
    if (reset) begin
      value <= 31'h0;
    end else if (_T_10) begin
      value <= 31'h0;
    end else begin
      value <= _T_12;
    end
    if (reset) begin
      q_data_sz <= 2'h3;
    end else begin
      q_data_sz <= _T_70;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_89) begin
          $fwrite(32'h80000002,"Assertion failed\n    at bridge.scala:168 assert ((~q_data_sz).orR =/= 0.U || !io.out.resp.valid)\n"); // @[bridge.scala 168:10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_89) begin
          $fatal; // @[bridge.scala 168:10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SimICache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input         io_in_req_bits_is_cached,
  input  [31:0] io_in_req_bits_addr,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [31:0] io_in_resp_bits_data,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output        io_out_req_bits_is_cached,
  output [31:0] io_out_req_bits_addr,
  output [1:0]  io_out_req_bits_len,
  output [3:0]  io_out_req_bits_strb,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [31:0] io_out_resp_bits_data,
  input         io_br_flush,
  input         io_ex_flush,
  input         io_control_valid,
  input  [2:0]  io_control_bits_op,
  input  [31:0] io_control_bits_addr
);
  reg  cache_v [0:255]; // @[icache.scala 91:18]
  reg [31:0] _RAND_0;
  wire  cache_v_s1_entry_r_data; // @[icache.scala 91:18]
  wire [7:0] cache_v_s1_entry_r_addr; // @[icache.scala 91:18]
  wire  cache_v__T_8_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_8_addr; // @[icache.scala 91:18]
  wire  cache_v__T_8_mask; // @[icache.scala 91:18]
  wire  cache_v__T_8_en; // @[icache.scala 91:18]
  wire  cache_v__T_10_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_10_addr; // @[icache.scala 91:18]
  wire  cache_v__T_10_mask; // @[icache.scala 91:18]
  wire  cache_v__T_10_en; // @[icache.scala 91:18]
  wire  cache_v__T_11_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_11_addr; // @[icache.scala 91:18]
  wire  cache_v__T_11_mask; // @[icache.scala 91:18]
  wire  cache_v__T_11_en; // @[icache.scala 91:18]
  wire  cache_v__T_12_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_12_addr; // @[icache.scala 91:18]
  wire  cache_v__T_12_mask; // @[icache.scala 91:18]
  wire  cache_v__T_12_en; // @[icache.scala 91:18]
  wire  cache_v__T_13_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_13_addr; // @[icache.scala 91:18]
  wire  cache_v__T_13_mask; // @[icache.scala 91:18]
  wire  cache_v__T_13_en; // @[icache.scala 91:18]
  wire  cache_v__T_14_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_14_addr; // @[icache.scala 91:18]
  wire  cache_v__T_14_mask; // @[icache.scala 91:18]
  wire  cache_v__T_14_en; // @[icache.scala 91:18]
  wire  cache_v__T_15_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_15_addr; // @[icache.scala 91:18]
  wire  cache_v__T_15_mask; // @[icache.scala 91:18]
  wire  cache_v__T_15_en; // @[icache.scala 91:18]
  wire  cache_v__T_16_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_16_addr; // @[icache.scala 91:18]
  wire  cache_v__T_16_mask; // @[icache.scala 91:18]
  wire  cache_v__T_16_en; // @[icache.scala 91:18]
  wire  cache_v__T_17_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_17_addr; // @[icache.scala 91:18]
  wire  cache_v__T_17_mask; // @[icache.scala 91:18]
  wire  cache_v__T_17_en; // @[icache.scala 91:18]
  wire  cache_v__T_18_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_18_addr; // @[icache.scala 91:18]
  wire  cache_v__T_18_mask; // @[icache.scala 91:18]
  wire  cache_v__T_18_en; // @[icache.scala 91:18]
  wire  cache_v__T_19_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_19_addr; // @[icache.scala 91:18]
  wire  cache_v__T_19_mask; // @[icache.scala 91:18]
  wire  cache_v__T_19_en; // @[icache.scala 91:18]
  wire  cache_v__T_20_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_20_addr; // @[icache.scala 91:18]
  wire  cache_v__T_20_mask; // @[icache.scala 91:18]
  wire  cache_v__T_20_en; // @[icache.scala 91:18]
  wire  cache_v__T_21_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_21_addr; // @[icache.scala 91:18]
  wire  cache_v__T_21_mask; // @[icache.scala 91:18]
  wire  cache_v__T_21_en; // @[icache.scala 91:18]
  wire  cache_v__T_22_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_22_addr; // @[icache.scala 91:18]
  wire  cache_v__T_22_mask; // @[icache.scala 91:18]
  wire  cache_v__T_22_en; // @[icache.scala 91:18]
  wire  cache_v__T_23_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_23_addr; // @[icache.scala 91:18]
  wire  cache_v__T_23_mask; // @[icache.scala 91:18]
  wire  cache_v__T_23_en; // @[icache.scala 91:18]
  wire  cache_v__T_24_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_24_addr; // @[icache.scala 91:18]
  wire  cache_v__T_24_mask; // @[icache.scala 91:18]
  wire  cache_v__T_24_en; // @[icache.scala 91:18]
  wire  cache_v__T_25_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_25_addr; // @[icache.scala 91:18]
  wire  cache_v__T_25_mask; // @[icache.scala 91:18]
  wire  cache_v__T_25_en; // @[icache.scala 91:18]
  wire  cache_v__T_26_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_26_addr; // @[icache.scala 91:18]
  wire  cache_v__T_26_mask; // @[icache.scala 91:18]
  wire  cache_v__T_26_en; // @[icache.scala 91:18]
  wire  cache_v__T_27_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_27_addr; // @[icache.scala 91:18]
  wire  cache_v__T_27_mask; // @[icache.scala 91:18]
  wire  cache_v__T_27_en; // @[icache.scala 91:18]
  wire  cache_v__T_28_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_28_addr; // @[icache.scala 91:18]
  wire  cache_v__T_28_mask; // @[icache.scala 91:18]
  wire  cache_v__T_28_en; // @[icache.scala 91:18]
  wire  cache_v__T_29_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_29_addr; // @[icache.scala 91:18]
  wire  cache_v__T_29_mask; // @[icache.scala 91:18]
  wire  cache_v__T_29_en; // @[icache.scala 91:18]
  wire  cache_v__T_30_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_30_addr; // @[icache.scala 91:18]
  wire  cache_v__T_30_mask; // @[icache.scala 91:18]
  wire  cache_v__T_30_en; // @[icache.scala 91:18]
  wire  cache_v__T_31_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_31_addr; // @[icache.scala 91:18]
  wire  cache_v__T_31_mask; // @[icache.scala 91:18]
  wire  cache_v__T_31_en; // @[icache.scala 91:18]
  wire  cache_v__T_32_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_32_addr; // @[icache.scala 91:18]
  wire  cache_v__T_32_mask; // @[icache.scala 91:18]
  wire  cache_v__T_32_en; // @[icache.scala 91:18]
  wire  cache_v__T_33_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_33_addr; // @[icache.scala 91:18]
  wire  cache_v__T_33_mask; // @[icache.scala 91:18]
  wire  cache_v__T_33_en; // @[icache.scala 91:18]
  wire  cache_v__T_34_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_34_addr; // @[icache.scala 91:18]
  wire  cache_v__T_34_mask; // @[icache.scala 91:18]
  wire  cache_v__T_34_en; // @[icache.scala 91:18]
  wire  cache_v__T_35_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_35_addr; // @[icache.scala 91:18]
  wire  cache_v__T_35_mask; // @[icache.scala 91:18]
  wire  cache_v__T_35_en; // @[icache.scala 91:18]
  wire  cache_v__T_36_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_36_addr; // @[icache.scala 91:18]
  wire  cache_v__T_36_mask; // @[icache.scala 91:18]
  wire  cache_v__T_36_en; // @[icache.scala 91:18]
  wire  cache_v__T_37_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_37_addr; // @[icache.scala 91:18]
  wire  cache_v__T_37_mask; // @[icache.scala 91:18]
  wire  cache_v__T_37_en; // @[icache.scala 91:18]
  wire  cache_v__T_38_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_38_addr; // @[icache.scala 91:18]
  wire  cache_v__T_38_mask; // @[icache.scala 91:18]
  wire  cache_v__T_38_en; // @[icache.scala 91:18]
  wire  cache_v__T_39_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_39_addr; // @[icache.scala 91:18]
  wire  cache_v__T_39_mask; // @[icache.scala 91:18]
  wire  cache_v__T_39_en; // @[icache.scala 91:18]
  wire  cache_v__T_40_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_40_addr; // @[icache.scala 91:18]
  wire  cache_v__T_40_mask; // @[icache.scala 91:18]
  wire  cache_v__T_40_en; // @[icache.scala 91:18]
  wire  cache_v__T_41_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_41_addr; // @[icache.scala 91:18]
  wire  cache_v__T_41_mask; // @[icache.scala 91:18]
  wire  cache_v__T_41_en; // @[icache.scala 91:18]
  wire  cache_v__T_42_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_42_addr; // @[icache.scala 91:18]
  wire  cache_v__T_42_mask; // @[icache.scala 91:18]
  wire  cache_v__T_42_en; // @[icache.scala 91:18]
  wire  cache_v__T_43_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_43_addr; // @[icache.scala 91:18]
  wire  cache_v__T_43_mask; // @[icache.scala 91:18]
  wire  cache_v__T_43_en; // @[icache.scala 91:18]
  wire  cache_v__T_44_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_44_addr; // @[icache.scala 91:18]
  wire  cache_v__T_44_mask; // @[icache.scala 91:18]
  wire  cache_v__T_44_en; // @[icache.scala 91:18]
  wire  cache_v__T_45_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_45_addr; // @[icache.scala 91:18]
  wire  cache_v__T_45_mask; // @[icache.scala 91:18]
  wire  cache_v__T_45_en; // @[icache.scala 91:18]
  wire  cache_v__T_46_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_46_addr; // @[icache.scala 91:18]
  wire  cache_v__T_46_mask; // @[icache.scala 91:18]
  wire  cache_v__T_46_en; // @[icache.scala 91:18]
  wire  cache_v__T_47_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_47_addr; // @[icache.scala 91:18]
  wire  cache_v__T_47_mask; // @[icache.scala 91:18]
  wire  cache_v__T_47_en; // @[icache.scala 91:18]
  wire  cache_v__T_48_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_48_addr; // @[icache.scala 91:18]
  wire  cache_v__T_48_mask; // @[icache.scala 91:18]
  wire  cache_v__T_48_en; // @[icache.scala 91:18]
  wire  cache_v__T_49_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_49_addr; // @[icache.scala 91:18]
  wire  cache_v__T_49_mask; // @[icache.scala 91:18]
  wire  cache_v__T_49_en; // @[icache.scala 91:18]
  wire  cache_v__T_50_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_50_addr; // @[icache.scala 91:18]
  wire  cache_v__T_50_mask; // @[icache.scala 91:18]
  wire  cache_v__T_50_en; // @[icache.scala 91:18]
  wire  cache_v__T_51_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_51_addr; // @[icache.scala 91:18]
  wire  cache_v__T_51_mask; // @[icache.scala 91:18]
  wire  cache_v__T_51_en; // @[icache.scala 91:18]
  wire  cache_v__T_52_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_52_addr; // @[icache.scala 91:18]
  wire  cache_v__T_52_mask; // @[icache.scala 91:18]
  wire  cache_v__T_52_en; // @[icache.scala 91:18]
  wire  cache_v__T_53_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_53_addr; // @[icache.scala 91:18]
  wire  cache_v__T_53_mask; // @[icache.scala 91:18]
  wire  cache_v__T_53_en; // @[icache.scala 91:18]
  wire  cache_v__T_54_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_54_addr; // @[icache.scala 91:18]
  wire  cache_v__T_54_mask; // @[icache.scala 91:18]
  wire  cache_v__T_54_en; // @[icache.scala 91:18]
  wire  cache_v__T_55_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_55_addr; // @[icache.scala 91:18]
  wire  cache_v__T_55_mask; // @[icache.scala 91:18]
  wire  cache_v__T_55_en; // @[icache.scala 91:18]
  wire  cache_v__T_56_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_56_addr; // @[icache.scala 91:18]
  wire  cache_v__T_56_mask; // @[icache.scala 91:18]
  wire  cache_v__T_56_en; // @[icache.scala 91:18]
  wire  cache_v__T_57_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_57_addr; // @[icache.scala 91:18]
  wire  cache_v__T_57_mask; // @[icache.scala 91:18]
  wire  cache_v__T_57_en; // @[icache.scala 91:18]
  wire  cache_v__T_58_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_58_addr; // @[icache.scala 91:18]
  wire  cache_v__T_58_mask; // @[icache.scala 91:18]
  wire  cache_v__T_58_en; // @[icache.scala 91:18]
  wire  cache_v__T_59_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_59_addr; // @[icache.scala 91:18]
  wire  cache_v__T_59_mask; // @[icache.scala 91:18]
  wire  cache_v__T_59_en; // @[icache.scala 91:18]
  wire  cache_v__T_60_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_60_addr; // @[icache.scala 91:18]
  wire  cache_v__T_60_mask; // @[icache.scala 91:18]
  wire  cache_v__T_60_en; // @[icache.scala 91:18]
  wire  cache_v__T_61_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_61_addr; // @[icache.scala 91:18]
  wire  cache_v__T_61_mask; // @[icache.scala 91:18]
  wire  cache_v__T_61_en; // @[icache.scala 91:18]
  wire  cache_v__T_62_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_62_addr; // @[icache.scala 91:18]
  wire  cache_v__T_62_mask; // @[icache.scala 91:18]
  wire  cache_v__T_62_en; // @[icache.scala 91:18]
  wire  cache_v__T_63_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_63_addr; // @[icache.scala 91:18]
  wire  cache_v__T_63_mask; // @[icache.scala 91:18]
  wire  cache_v__T_63_en; // @[icache.scala 91:18]
  wire  cache_v__T_64_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_64_addr; // @[icache.scala 91:18]
  wire  cache_v__T_64_mask; // @[icache.scala 91:18]
  wire  cache_v__T_64_en; // @[icache.scala 91:18]
  wire  cache_v__T_65_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_65_addr; // @[icache.scala 91:18]
  wire  cache_v__T_65_mask; // @[icache.scala 91:18]
  wire  cache_v__T_65_en; // @[icache.scala 91:18]
  wire  cache_v__T_66_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_66_addr; // @[icache.scala 91:18]
  wire  cache_v__T_66_mask; // @[icache.scala 91:18]
  wire  cache_v__T_66_en; // @[icache.scala 91:18]
  wire  cache_v__T_67_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_67_addr; // @[icache.scala 91:18]
  wire  cache_v__T_67_mask; // @[icache.scala 91:18]
  wire  cache_v__T_67_en; // @[icache.scala 91:18]
  wire  cache_v__T_68_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_68_addr; // @[icache.scala 91:18]
  wire  cache_v__T_68_mask; // @[icache.scala 91:18]
  wire  cache_v__T_68_en; // @[icache.scala 91:18]
  wire  cache_v__T_69_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_69_addr; // @[icache.scala 91:18]
  wire  cache_v__T_69_mask; // @[icache.scala 91:18]
  wire  cache_v__T_69_en; // @[icache.scala 91:18]
  wire  cache_v__T_70_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_70_addr; // @[icache.scala 91:18]
  wire  cache_v__T_70_mask; // @[icache.scala 91:18]
  wire  cache_v__T_70_en; // @[icache.scala 91:18]
  wire  cache_v__T_71_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_71_addr; // @[icache.scala 91:18]
  wire  cache_v__T_71_mask; // @[icache.scala 91:18]
  wire  cache_v__T_71_en; // @[icache.scala 91:18]
  wire  cache_v__T_72_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_72_addr; // @[icache.scala 91:18]
  wire  cache_v__T_72_mask; // @[icache.scala 91:18]
  wire  cache_v__T_72_en; // @[icache.scala 91:18]
  wire  cache_v__T_73_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_73_addr; // @[icache.scala 91:18]
  wire  cache_v__T_73_mask; // @[icache.scala 91:18]
  wire  cache_v__T_73_en; // @[icache.scala 91:18]
  wire  cache_v__T_74_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_74_addr; // @[icache.scala 91:18]
  wire  cache_v__T_74_mask; // @[icache.scala 91:18]
  wire  cache_v__T_74_en; // @[icache.scala 91:18]
  wire  cache_v__T_75_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_75_addr; // @[icache.scala 91:18]
  wire  cache_v__T_75_mask; // @[icache.scala 91:18]
  wire  cache_v__T_75_en; // @[icache.scala 91:18]
  wire  cache_v__T_76_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_76_addr; // @[icache.scala 91:18]
  wire  cache_v__T_76_mask; // @[icache.scala 91:18]
  wire  cache_v__T_76_en; // @[icache.scala 91:18]
  wire  cache_v__T_77_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_77_addr; // @[icache.scala 91:18]
  wire  cache_v__T_77_mask; // @[icache.scala 91:18]
  wire  cache_v__T_77_en; // @[icache.scala 91:18]
  wire  cache_v__T_78_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_78_addr; // @[icache.scala 91:18]
  wire  cache_v__T_78_mask; // @[icache.scala 91:18]
  wire  cache_v__T_78_en; // @[icache.scala 91:18]
  wire  cache_v__T_79_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_79_addr; // @[icache.scala 91:18]
  wire  cache_v__T_79_mask; // @[icache.scala 91:18]
  wire  cache_v__T_79_en; // @[icache.scala 91:18]
  wire  cache_v__T_80_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_80_addr; // @[icache.scala 91:18]
  wire  cache_v__T_80_mask; // @[icache.scala 91:18]
  wire  cache_v__T_80_en; // @[icache.scala 91:18]
  wire  cache_v__T_81_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_81_addr; // @[icache.scala 91:18]
  wire  cache_v__T_81_mask; // @[icache.scala 91:18]
  wire  cache_v__T_81_en; // @[icache.scala 91:18]
  wire  cache_v__T_82_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_82_addr; // @[icache.scala 91:18]
  wire  cache_v__T_82_mask; // @[icache.scala 91:18]
  wire  cache_v__T_82_en; // @[icache.scala 91:18]
  wire  cache_v__T_83_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_83_addr; // @[icache.scala 91:18]
  wire  cache_v__T_83_mask; // @[icache.scala 91:18]
  wire  cache_v__T_83_en; // @[icache.scala 91:18]
  wire  cache_v__T_84_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_84_addr; // @[icache.scala 91:18]
  wire  cache_v__T_84_mask; // @[icache.scala 91:18]
  wire  cache_v__T_84_en; // @[icache.scala 91:18]
  wire  cache_v__T_85_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_85_addr; // @[icache.scala 91:18]
  wire  cache_v__T_85_mask; // @[icache.scala 91:18]
  wire  cache_v__T_85_en; // @[icache.scala 91:18]
  wire  cache_v__T_86_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_86_addr; // @[icache.scala 91:18]
  wire  cache_v__T_86_mask; // @[icache.scala 91:18]
  wire  cache_v__T_86_en; // @[icache.scala 91:18]
  wire  cache_v__T_87_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_87_addr; // @[icache.scala 91:18]
  wire  cache_v__T_87_mask; // @[icache.scala 91:18]
  wire  cache_v__T_87_en; // @[icache.scala 91:18]
  wire  cache_v__T_88_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_88_addr; // @[icache.scala 91:18]
  wire  cache_v__T_88_mask; // @[icache.scala 91:18]
  wire  cache_v__T_88_en; // @[icache.scala 91:18]
  wire  cache_v__T_89_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_89_addr; // @[icache.scala 91:18]
  wire  cache_v__T_89_mask; // @[icache.scala 91:18]
  wire  cache_v__T_89_en; // @[icache.scala 91:18]
  wire  cache_v__T_90_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_90_addr; // @[icache.scala 91:18]
  wire  cache_v__T_90_mask; // @[icache.scala 91:18]
  wire  cache_v__T_90_en; // @[icache.scala 91:18]
  wire  cache_v__T_91_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_91_addr; // @[icache.scala 91:18]
  wire  cache_v__T_91_mask; // @[icache.scala 91:18]
  wire  cache_v__T_91_en; // @[icache.scala 91:18]
  wire  cache_v__T_92_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_92_addr; // @[icache.scala 91:18]
  wire  cache_v__T_92_mask; // @[icache.scala 91:18]
  wire  cache_v__T_92_en; // @[icache.scala 91:18]
  wire  cache_v__T_93_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_93_addr; // @[icache.scala 91:18]
  wire  cache_v__T_93_mask; // @[icache.scala 91:18]
  wire  cache_v__T_93_en; // @[icache.scala 91:18]
  wire  cache_v__T_94_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_94_addr; // @[icache.scala 91:18]
  wire  cache_v__T_94_mask; // @[icache.scala 91:18]
  wire  cache_v__T_94_en; // @[icache.scala 91:18]
  wire  cache_v__T_95_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_95_addr; // @[icache.scala 91:18]
  wire  cache_v__T_95_mask; // @[icache.scala 91:18]
  wire  cache_v__T_95_en; // @[icache.scala 91:18]
  wire  cache_v__T_96_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_96_addr; // @[icache.scala 91:18]
  wire  cache_v__T_96_mask; // @[icache.scala 91:18]
  wire  cache_v__T_96_en; // @[icache.scala 91:18]
  wire  cache_v__T_97_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_97_addr; // @[icache.scala 91:18]
  wire  cache_v__T_97_mask; // @[icache.scala 91:18]
  wire  cache_v__T_97_en; // @[icache.scala 91:18]
  wire  cache_v__T_98_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_98_addr; // @[icache.scala 91:18]
  wire  cache_v__T_98_mask; // @[icache.scala 91:18]
  wire  cache_v__T_98_en; // @[icache.scala 91:18]
  wire  cache_v__T_99_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_99_addr; // @[icache.scala 91:18]
  wire  cache_v__T_99_mask; // @[icache.scala 91:18]
  wire  cache_v__T_99_en; // @[icache.scala 91:18]
  wire  cache_v__T_100_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_100_addr; // @[icache.scala 91:18]
  wire  cache_v__T_100_mask; // @[icache.scala 91:18]
  wire  cache_v__T_100_en; // @[icache.scala 91:18]
  wire  cache_v__T_101_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_101_addr; // @[icache.scala 91:18]
  wire  cache_v__T_101_mask; // @[icache.scala 91:18]
  wire  cache_v__T_101_en; // @[icache.scala 91:18]
  wire  cache_v__T_102_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_102_addr; // @[icache.scala 91:18]
  wire  cache_v__T_102_mask; // @[icache.scala 91:18]
  wire  cache_v__T_102_en; // @[icache.scala 91:18]
  wire  cache_v__T_103_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_103_addr; // @[icache.scala 91:18]
  wire  cache_v__T_103_mask; // @[icache.scala 91:18]
  wire  cache_v__T_103_en; // @[icache.scala 91:18]
  wire  cache_v__T_104_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_104_addr; // @[icache.scala 91:18]
  wire  cache_v__T_104_mask; // @[icache.scala 91:18]
  wire  cache_v__T_104_en; // @[icache.scala 91:18]
  wire  cache_v__T_105_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_105_addr; // @[icache.scala 91:18]
  wire  cache_v__T_105_mask; // @[icache.scala 91:18]
  wire  cache_v__T_105_en; // @[icache.scala 91:18]
  wire  cache_v__T_106_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_106_addr; // @[icache.scala 91:18]
  wire  cache_v__T_106_mask; // @[icache.scala 91:18]
  wire  cache_v__T_106_en; // @[icache.scala 91:18]
  wire  cache_v__T_107_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_107_addr; // @[icache.scala 91:18]
  wire  cache_v__T_107_mask; // @[icache.scala 91:18]
  wire  cache_v__T_107_en; // @[icache.scala 91:18]
  wire  cache_v__T_108_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_108_addr; // @[icache.scala 91:18]
  wire  cache_v__T_108_mask; // @[icache.scala 91:18]
  wire  cache_v__T_108_en; // @[icache.scala 91:18]
  wire  cache_v__T_109_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_109_addr; // @[icache.scala 91:18]
  wire  cache_v__T_109_mask; // @[icache.scala 91:18]
  wire  cache_v__T_109_en; // @[icache.scala 91:18]
  wire  cache_v__T_110_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_110_addr; // @[icache.scala 91:18]
  wire  cache_v__T_110_mask; // @[icache.scala 91:18]
  wire  cache_v__T_110_en; // @[icache.scala 91:18]
  wire  cache_v__T_111_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_111_addr; // @[icache.scala 91:18]
  wire  cache_v__T_111_mask; // @[icache.scala 91:18]
  wire  cache_v__T_111_en; // @[icache.scala 91:18]
  wire  cache_v__T_112_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_112_addr; // @[icache.scala 91:18]
  wire  cache_v__T_112_mask; // @[icache.scala 91:18]
  wire  cache_v__T_112_en; // @[icache.scala 91:18]
  wire  cache_v__T_113_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_113_addr; // @[icache.scala 91:18]
  wire  cache_v__T_113_mask; // @[icache.scala 91:18]
  wire  cache_v__T_113_en; // @[icache.scala 91:18]
  wire  cache_v__T_114_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_114_addr; // @[icache.scala 91:18]
  wire  cache_v__T_114_mask; // @[icache.scala 91:18]
  wire  cache_v__T_114_en; // @[icache.scala 91:18]
  wire  cache_v__T_115_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_115_addr; // @[icache.scala 91:18]
  wire  cache_v__T_115_mask; // @[icache.scala 91:18]
  wire  cache_v__T_115_en; // @[icache.scala 91:18]
  wire  cache_v__T_116_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_116_addr; // @[icache.scala 91:18]
  wire  cache_v__T_116_mask; // @[icache.scala 91:18]
  wire  cache_v__T_116_en; // @[icache.scala 91:18]
  wire  cache_v__T_117_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_117_addr; // @[icache.scala 91:18]
  wire  cache_v__T_117_mask; // @[icache.scala 91:18]
  wire  cache_v__T_117_en; // @[icache.scala 91:18]
  wire  cache_v__T_118_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_118_addr; // @[icache.scala 91:18]
  wire  cache_v__T_118_mask; // @[icache.scala 91:18]
  wire  cache_v__T_118_en; // @[icache.scala 91:18]
  wire  cache_v__T_119_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_119_addr; // @[icache.scala 91:18]
  wire  cache_v__T_119_mask; // @[icache.scala 91:18]
  wire  cache_v__T_119_en; // @[icache.scala 91:18]
  wire  cache_v__T_120_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_120_addr; // @[icache.scala 91:18]
  wire  cache_v__T_120_mask; // @[icache.scala 91:18]
  wire  cache_v__T_120_en; // @[icache.scala 91:18]
  wire  cache_v__T_121_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_121_addr; // @[icache.scala 91:18]
  wire  cache_v__T_121_mask; // @[icache.scala 91:18]
  wire  cache_v__T_121_en; // @[icache.scala 91:18]
  wire  cache_v__T_122_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_122_addr; // @[icache.scala 91:18]
  wire  cache_v__T_122_mask; // @[icache.scala 91:18]
  wire  cache_v__T_122_en; // @[icache.scala 91:18]
  wire  cache_v__T_123_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_123_addr; // @[icache.scala 91:18]
  wire  cache_v__T_123_mask; // @[icache.scala 91:18]
  wire  cache_v__T_123_en; // @[icache.scala 91:18]
  wire  cache_v__T_124_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_124_addr; // @[icache.scala 91:18]
  wire  cache_v__T_124_mask; // @[icache.scala 91:18]
  wire  cache_v__T_124_en; // @[icache.scala 91:18]
  wire  cache_v__T_125_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_125_addr; // @[icache.scala 91:18]
  wire  cache_v__T_125_mask; // @[icache.scala 91:18]
  wire  cache_v__T_125_en; // @[icache.scala 91:18]
  wire  cache_v__T_126_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_126_addr; // @[icache.scala 91:18]
  wire  cache_v__T_126_mask; // @[icache.scala 91:18]
  wire  cache_v__T_126_en; // @[icache.scala 91:18]
  wire  cache_v__T_127_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_127_addr; // @[icache.scala 91:18]
  wire  cache_v__T_127_mask; // @[icache.scala 91:18]
  wire  cache_v__T_127_en; // @[icache.scala 91:18]
  wire  cache_v__T_128_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_128_addr; // @[icache.scala 91:18]
  wire  cache_v__T_128_mask; // @[icache.scala 91:18]
  wire  cache_v__T_128_en; // @[icache.scala 91:18]
  wire  cache_v__T_129_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_129_addr; // @[icache.scala 91:18]
  wire  cache_v__T_129_mask; // @[icache.scala 91:18]
  wire  cache_v__T_129_en; // @[icache.scala 91:18]
  wire  cache_v__T_130_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_130_addr; // @[icache.scala 91:18]
  wire  cache_v__T_130_mask; // @[icache.scala 91:18]
  wire  cache_v__T_130_en; // @[icache.scala 91:18]
  wire  cache_v__T_131_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_131_addr; // @[icache.scala 91:18]
  wire  cache_v__T_131_mask; // @[icache.scala 91:18]
  wire  cache_v__T_131_en; // @[icache.scala 91:18]
  wire  cache_v__T_132_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_132_addr; // @[icache.scala 91:18]
  wire  cache_v__T_132_mask; // @[icache.scala 91:18]
  wire  cache_v__T_132_en; // @[icache.scala 91:18]
  wire  cache_v__T_133_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_133_addr; // @[icache.scala 91:18]
  wire  cache_v__T_133_mask; // @[icache.scala 91:18]
  wire  cache_v__T_133_en; // @[icache.scala 91:18]
  wire  cache_v__T_134_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_134_addr; // @[icache.scala 91:18]
  wire  cache_v__T_134_mask; // @[icache.scala 91:18]
  wire  cache_v__T_134_en; // @[icache.scala 91:18]
  wire  cache_v__T_135_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_135_addr; // @[icache.scala 91:18]
  wire  cache_v__T_135_mask; // @[icache.scala 91:18]
  wire  cache_v__T_135_en; // @[icache.scala 91:18]
  wire  cache_v__T_136_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_136_addr; // @[icache.scala 91:18]
  wire  cache_v__T_136_mask; // @[icache.scala 91:18]
  wire  cache_v__T_136_en; // @[icache.scala 91:18]
  wire  cache_v__T_137_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_137_addr; // @[icache.scala 91:18]
  wire  cache_v__T_137_mask; // @[icache.scala 91:18]
  wire  cache_v__T_137_en; // @[icache.scala 91:18]
  wire  cache_v__T_138_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_138_addr; // @[icache.scala 91:18]
  wire  cache_v__T_138_mask; // @[icache.scala 91:18]
  wire  cache_v__T_138_en; // @[icache.scala 91:18]
  wire  cache_v__T_139_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_139_addr; // @[icache.scala 91:18]
  wire  cache_v__T_139_mask; // @[icache.scala 91:18]
  wire  cache_v__T_139_en; // @[icache.scala 91:18]
  wire  cache_v__T_140_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_140_addr; // @[icache.scala 91:18]
  wire  cache_v__T_140_mask; // @[icache.scala 91:18]
  wire  cache_v__T_140_en; // @[icache.scala 91:18]
  wire  cache_v__T_141_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_141_addr; // @[icache.scala 91:18]
  wire  cache_v__T_141_mask; // @[icache.scala 91:18]
  wire  cache_v__T_141_en; // @[icache.scala 91:18]
  wire  cache_v__T_142_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_142_addr; // @[icache.scala 91:18]
  wire  cache_v__T_142_mask; // @[icache.scala 91:18]
  wire  cache_v__T_142_en; // @[icache.scala 91:18]
  wire  cache_v__T_143_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_143_addr; // @[icache.scala 91:18]
  wire  cache_v__T_143_mask; // @[icache.scala 91:18]
  wire  cache_v__T_143_en; // @[icache.scala 91:18]
  wire  cache_v__T_144_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_144_addr; // @[icache.scala 91:18]
  wire  cache_v__T_144_mask; // @[icache.scala 91:18]
  wire  cache_v__T_144_en; // @[icache.scala 91:18]
  wire  cache_v__T_145_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_145_addr; // @[icache.scala 91:18]
  wire  cache_v__T_145_mask; // @[icache.scala 91:18]
  wire  cache_v__T_145_en; // @[icache.scala 91:18]
  wire  cache_v__T_146_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_146_addr; // @[icache.scala 91:18]
  wire  cache_v__T_146_mask; // @[icache.scala 91:18]
  wire  cache_v__T_146_en; // @[icache.scala 91:18]
  wire  cache_v__T_147_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_147_addr; // @[icache.scala 91:18]
  wire  cache_v__T_147_mask; // @[icache.scala 91:18]
  wire  cache_v__T_147_en; // @[icache.scala 91:18]
  wire  cache_v__T_148_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_148_addr; // @[icache.scala 91:18]
  wire  cache_v__T_148_mask; // @[icache.scala 91:18]
  wire  cache_v__T_148_en; // @[icache.scala 91:18]
  wire  cache_v__T_149_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_149_addr; // @[icache.scala 91:18]
  wire  cache_v__T_149_mask; // @[icache.scala 91:18]
  wire  cache_v__T_149_en; // @[icache.scala 91:18]
  wire  cache_v__T_150_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_150_addr; // @[icache.scala 91:18]
  wire  cache_v__T_150_mask; // @[icache.scala 91:18]
  wire  cache_v__T_150_en; // @[icache.scala 91:18]
  wire  cache_v__T_151_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_151_addr; // @[icache.scala 91:18]
  wire  cache_v__T_151_mask; // @[icache.scala 91:18]
  wire  cache_v__T_151_en; // @[icache.scala 91:18]
  wire  cache_v__T_152_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_152_addr; // @[icache.scala 91:18]
  wire  cache_v__T_152_mask; // @[icache.scala 91:18]
  wire  cache_v__T_152_en; // @[icache.scala 91:18]
  wire  cache_v__T_153_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_153_addr; // @[icache.scala 91:18]
  wire  cache_v__T_153_mask; // @[icache.scala 91:18]
  wire  cache_v__T_153_en; // @[icache.scala 91:18]
  wire  cache_v__T_154_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_154_addr; // @[icache.scala 91:18]
  wire  cache_v__T_154_mask; // @[icache.scala 91:18]
  wire  cache_v__T_154_en; // @[icache.scala 91:18]
  wire  cache_v__T_155_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_155_addr; // @[icache.scala 91:18]
  wire  cache_v__T_155_mask; // @[icache.scala 91:18]
  wire  cache_v__T_155_en; // @[icache.scala 91:18]
  wire  cache_v__T_156_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_156_addr; // @[icache.scala 91:18]
  wire  cache_v__T_156_mask; // @[icache.scala 91:18]
  wire  cache_v__T_156_en; // @[icache.scala 91:18]
  wire  cache_v__T_157_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_157_addr; // @[icache.scala 91:18]
  wire  cache_v__T_157_mask; // @[icache.scala 91:18]
  wire  cache_v__T_157_en; // @[icache.scala 91:18]
  wire  cache_v__T_158_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_158_addr; // @[icache.scala 91:18]
  wire  cache_v__T_158_mask; // @[icache.scala 91:18]
  wire  cache_v__T_158_en; // @[icache.scala 91:18]
  wire  cache_v__T_159_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_159_addr; // @[icache.scala 91:18]
  wire  cache_v__T_159_mask; // @[icache.scala 91:18]
  wire  cache_v__T_159_en; // @[icache.scala 91:18]
  wire  cache_v__T_160_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_160_addr; // @[icache.scala 91:18]
  wire  cache_v__T_160_mask; // @[icache.scala 91:18]
  wire  cache_v__T_160_en; // @[icache.scala 91:18]
  wire  cache_v__T_161_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_161_addr; // @[icache.scala 91:18]
  wire  cache_v__T_161_mask; // @[icache.scala 91:18]
  wire  cache_v__T_161_en; // @[icache.scala 91:18]
  wire  cache_v__T_162_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_162_addr; // @[icache.scala 91:18]
  wire  cache_v__T_162_mask; // @[icache.scala 91:18]
  wire  cache_v__T_162_en; // @[icache.scala 91:18]
  wire  cache_v__T_163_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_163_addr; // @[icache.scala 91:18]
  wire  cache_v__T_163_mask; // @[icache.scala 91:18]
  wire  cache_v__T_163_en; // @[icache.scala 91:18]
  wire  cache_v__T_164_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_164_addr; // @[icache.scala 91:18]
  wire  cache_v__T_164_mask; // @[icache.scala 91:18]
  wire  cache_v__T_164_en; // @[icache.scala 91:18]
  wire  cache_v__T_165_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_165_addr; // @[icache.scala 91:18]
  wire  cache_v__T_165_mask; // @[icache.scala 91:18]
  wire  cache_v__T_165_en; // @[icache.scala 91:18]
  wire  cache_v__T_166_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_166_addr; // @[icache.scala 91:18]
  wire  cache_v__T_166_mask; // @[icache.scala 91:18]
  wire  cache_v__T_166_en; // @[icache.scala 91:18]
  wire  cache_v__T_167_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_167_addr; // @[icache.scala 91:18]
  wire  cache_v__T_167_mask; // @[icache.scala 91:18]
  wire  cache_v__T_167_en; // @[icache.scala 91:18]
  wire  cache_v__T_168_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_168_addr; // @[icache.scala 91:18]
  wire  cache_v__T_168_mask; // @[icache.scala 91:18]
  wire  cache_v__T_168_en; // @[icache.scala 91:18]
  wire  cache_v__T_169_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_169_addr; // @[icache.scala 91:18]
  wire  cache_v__T_169_mask; // @[icache.scala 91:18]
  wire  cache_v__T_169_en; // @[icache.scala 91:18]
  wire  cache_v__T_170_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_170_addr; // @[icache.scala 91:18]
  wire  cache_v__T_170_mask; // @[icache.scala 91:18]
  wire  cache_v__T_170_en; // @[icache.scala 91:18]
  wire  cache_v__T_171_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_171_addr; // @[icache.scala 91:18]
  wire  cache_v__T_171_mask; // @[icache.scala 91:18]
  wire  cache_v__T_171_en; // @[icache.scala 91:18]
  wire  cache_v__T_172_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_172_addr; // @[icache.scala 91:18]
  wire  cache_v__T_172_mask; // @[icache.scala 91:18]
  wire  cache_v__T_172_en; // @[icache.scala 91:18]
  wire  cache_v__T_173_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_173_addr; // @[icache.scala 91:18]
  wire  cache_v__T_173_mask; // @[icache.scala 91:18]
  wire  cache_v__T_173_en; // @[icache.scala 91:18]
  wire  cache_v__T_174_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_174_addr; // @[icache.scala 91:18]
  wire  cache_v__T_174_mask; // @[icache.scala 91:18]
  wire  cache_v__T_174_en; // @[icache.scala 91:18]
  wire  cache_v__T_175_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_175_addr; // @[icache.scala 91:18]
  wire  cache_v__T_175_mask; // @[icache.scala 91:18]
  wire  cache_v__T_175_en; // @[icache.scala 91:18]
  wire  cache_v__T_176_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_176_addr; // @[icache.scala 91:18]
  wire  cache_v__T_176_mask; // @[icache.scala 91:18]
  wire  cache_v__T_176_en; // @[icache.scala 91:18]
  wire  cache_v__T_177_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_177_addr; // @[icache.scala 91:18]
  wire  cache_v__T_177_mask; // @[icache.scala 91:18]
  wire  cache_v__T_177_en; // @[icache.scala 91:18]
  wire  cache_v__T_178_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_178_addr; // @[icache.scala 91:18]
  wire  cache_v__T_178_mask; // @[icache.scala 91:18]
  wire  cache_v__T_178_en; // @[icache.scala 91:18]
  wire  cache_v__T_179_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_179_addr; // @[icache.scala 91:18]
  wire  cache_v__T_179_mask; // @[icache.scala 91:18]
  wire  cache_v__T_179_en; // @[icache.scala 91:18]
  wire  cache_v__T_180_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_180_addr; // @[icache.scala 91:18]
  wire  cache_v__T_180_mask; // @[icache.scala 91:18]
  wire  cache_v__T_180_en; // @[icache.scala 91:18]
  wire  cache_v__T_181_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_181_addr; // @[icache.scala 91:18]
  wire  cache_v__T_181_mask; // @[icache.scala 91:18]
  wire  cache_v__T_181_en; // @[icache.scala 91:18]
  wire  cache_v__T_182_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_182_addr; // @[icache.scala 91:18]
  wire  cache_v__T_182_mask; // @[icache.scala 91:18]
  wire  cache_v__T_182_en; // @[icache.scala 91:18]
  wire  cache_v__T_183_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_183_addr; // @[icache.scala 91:18]
  wire  cache_v__T_183_mask; // @[icache.scala 91:18]
  wire  cache_v__T_183_en; // @[icache.scala 91:18]
  wire  cache_v__T_184_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_184_addr; // @[icache.scala 91:18]
  wire  cache_v__T_184_mask; // @[icache.scala 91:18]
  wire  cache_v__T_184_en; // @[icache.scala 91:18]
  wire  cache_v__T_185_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_185_addr; // @[icache.scala 91:18]
  wire  cache_v__T_185_mask; // @[icache.scala 91:18]
  wire  cache_v__T_185_en; // @[icache.scala 91:18]
  wire  cache_v__T_186_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_186_addr; // @[icache.scala 91:18]
  wire  cache_v__T_186_mask; // @[icache.scala 91:18]
  wire  cache_v__T_186_en; // @[icache.scala 91:18]
  wire  cache_v__T_187_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_187_addr; // @[icache.scala 91:18]
  wire  cache_v__T_187_mask; // @[icache.scala 91:18]
  wire  cache_v__T_187_en; // @[icache.scala 91:18]
  wire  cache_v__T_188_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_188_addr; // @[icache.scala 91:18]
  wire  cache_v__T_188_mask; // @[icache.scala 91:18]
  wire  cache_v__T_188_en; // @[icache.scala 91:18]
  wire  cache_v__T_189_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_189_addr; // @[icache.scala 91:18]
  wire  cache_v__T_189_mask; // @[icache.scala 91:18]
  wire  cache_v__T_189_en; // @[icache.scala 91:18]
  wire  cache_v__T_190_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_190_addr; // @[icache.scala 91:18]
  wire  cache_v__T_190_mask; // @[icache.scala 91:18]
  wire  cache_v__T_190_en; // @[icache.scala 91:18]
  wire  cache_v__T_191_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_191_addr; // @[icache.scala 91:18]
  wire  cache_v__T_191_mask; // @[icache.scala 91:18]
  wire  cache_v__T_191_en; // @[icache.scala 91:18]
  wire  cache_v__T_192_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_192_addr; // @[icache.scala 91:18]
  wire  cache_v__T_192_mask; // @[icache.scala 91:18]
  wire  cache_v__T_192_en; // @[icache.scala 91:18]
  wire  cache_v__T_193_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_193_addr; // @[icache.scala 91:18]
  wire  cache_v__T_193_mask; // @[icache.scala 91:18]
  wire  cache_v__T_193_en; // @[icache.scala 91:18]
  wire  cache_v__T_194_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_194_addr; // @[icache.scala 91:18]
  wire  cache_v__T_194_mask; // @[icache.scala 91:18]
  wire  cache_v__T_194_en; // @[icache.scala 91:18]
  wire  cache_v__T_195_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_195_addr; // @[icache.scala 91:18]
  wire  cache_v__T_195_mask; // @[icache.scala 91:18]
  wire  cache_v__T_195_en; // @[icache.scala 91:18]
  wire  cache_v__T_196_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_196_addr; // @[icache.scala 91:18]
  wire  cache_v__T_196_mask; // @[icache.scala 91:18]
  wire  cache_v__T_196_en; // @[icache.scala 91:18]
  wire  cache_v__T_197_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_197_addr; // @[icache.scala 91:18]
  wire  cache_v__T_197_mask; // @[icache.scala 91:18]
  wire  cache_v__T_197_en; // @[icache.scala 91:18]
  wire  cache_v__T_198_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_198_addr; // @[icache.scala 91:18]
  wire  cache_v__T_198_mask; // @[icache.scala 91:18]
  wire  cache_v__T_198_en; // @[icache.scala 91:18]
  wire  cache_v__T_199_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_199_addr; // @[icache.scala 91:18]
  wire  cache_v__T_199_mask; // @[icache.scala 91:18]
  wire  cache_v__T_199_en; // @[icache.scala 91:18]
  wire  cache_v__T_200_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_200_addr; // @[icache.scala 91:18]
  wire  cache_v__T_200_mask; // @[icache.scala 91:18]
  wire  cache_v__T_200_en; // @[icache.scala 91:18]
  wire  cache_v__T_201_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_201_addr; // @[icache.scala 91:18]
  wire  cache_v__T_201_mask; // @[icache.scala 91:18]
  wire  cache_v__T_201_en; // @[icache.scala 91:18]
  wire  cache_v__T_202_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_202_addr; // @[icache.scala 91:18]
  wire  cache_v__T_202_mask; // @[icache.scala 91:18]
  wire  cache_v__T_202_en; // @[icache.scala 91:18]
  wire  cache_v__T_203_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_203_addr; // @[icache.scala 91:18]
  wire  cache_v__T_203_mask; // @[icache.scala 91:18]
  wire  cache_v__T_203_en; // @[icache.scala 91:18]
  wire  cache_v__T_204_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_204_addr; // @[icache.scala 91:18]
  wire  cache_v__T_204_mask; // @[icache.scala 91:18]
  wire  cache_v__T_204_en; // @[icache.scala 91:18]
  wire  cache_v__T_205_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_205_addr; // @[icache.scala 91:18]
  wire  cache_v__T_205_mask; // @[icache.scala 91:18]
  wire  cache_v__T_205_en; // @[icache.scala 91:18]
  wire  cache_v__T_206_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_206_addr; // @[icache.scala 91:18]
  wire  cache_v__T_206_mask; // @[icache.scala 91:18]
  wire  cache_v__T_206_en; // @[icache.scala 91:18]
  wire  cache_v__T_207_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_207_addr; // @[icache.scala 91:18]
  wire  cache_v__T_207_mask; // @[icache.scala 91:18]
  wire  cache_v__T_207_en; // @[icache.scala 91:18]
  wire  cache_v__T_208_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_208_addr; // @[icache.scala 91:18]
  wire  cache_v__T_208_mask; // @[icache.scala 91:18]
  wire  cache_v__T_208_en; // @[icache.scala 91:18]
  wire  cache_v__T_209_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_209_addr; // @[icache.scala 91:18]
  wire  cache_v__T_209_mask; // @[icache.scala 91:18]
  wire  cache_v__T_209_en; // @[icache.scala 91:18]
  wire  cache_v__T_210_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_210_addr; // @[icache.scala 91:18]
  wire  cache_v__T_210_mask; // @[icache.scala 91:18]
  wire  cache_v__T_210_en; // @[icache.scala 91:18]
  wire  cache_v__T_211_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_211_addr; // @[icache.scala 91:18]
  wire  cache_v__T_211_mask; // @[icache.scala 91:18]
  wire  cache_v__T_211_en; // @[icache.scala 91:18]
  wire  cache_v__T_212_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_212_addr; // @[icache.scala 91:18]
  wire  cache_v__T_212_mask; // @[icache.scala 91:18]
  wire  cache_v__T_212_en; // @[icache.scala 91:18]
  wire  cache_v__T_213_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_213_addr; // @[icache.scala 91:18]
  wire  cache_v__T_213_mask; // @[icache.scala 91:18]
  wire  cache_v__T_213_en; // @[icache.scala 91:18]
  wire  cache_v__T_214_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_214_addr; // @[icache.scala 91:18]
  wire  cache_v__T_214_mask; // @[icache.scala 91:18]
  wire  cache_v__T_214_en; // @[icache.scala 91:18]
  wire  cache_v__T_215_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_215_addr; // @[icache.scala 91:18]
  wire  cache_v__T_215_mask; // @[icache.scala 91:18]
  wire  cache_v__T_215_en; // @[icache.scala 91:18]
  wire  cache_v__T_216_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_216_addr; // @[icache.scala 91:18]
  wire  cache_v__T_216_mask; // @[icache.scala 91:18]
  wire  cache_v__T_216_en; // @[icache.scala 91:18]
  wire  cache_v__T_217_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_217_addr; // @[icache.scala 91:18]
  wire  cache_v__T_217_mask; // @[icache.scala 91:18]
  wire  cache_v__T_217_en; // @[icache.scala 91:18]
  wire  cache_v__T_218_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_218_addr; // @[icache.scala 91:18]
  wire  cache_v__T_218_mask; // @[icache.scala 91:18]
  wire  cache_v__T_218_en; // @[icache.scala 91:18]
  wire  cache_v__T_219_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_219_addr; // @[icache.scala 91:18]
  wire  cache_v__T_219_mask; // @[icache.scala 91:18]
  wire  cache_v__T_219_en; // @[icache.scala 91:18]
  wire  cache_v__T_220_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_220_addr; // @[icache.scala 91:18]
  wire  cache_v__T_220_mask; // @[icache.scala 91:18]
  wire  cache_v__T_220_en; // @[icache.scala 91:18]
  wire  cache_v__T_221_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_221_addr; // @[icache.scala 91:18]
  wire  cache_v__T_221_mask; // @[icache.scala 91:18]
  wire  cache_v__T_221_en; // @[icache.scala 91:18]
  wire  cache_v__T_222_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_222_addr; // @[icache.scala 91:18]
  wire  cache_v__T_222_mask; // @[icache.scala 91:18]
  wire  cache_v__T_222_en; // @[icache.scala 91:18]
  wire  cache_v__T_223_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_223_addr; // @[icache.scala 91:18]
  wire  cache_v__T_223_mask; // @[icache.scala 91:18]
  wire  cache_v__T_223_en; // @[icache.scala 91:18]
  wire  cache_v__T_224_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_224_addr; // @[icache.scala 91:18]
  wire  cache_v__T_224_mask; // @[icache.scala 91:18]
  wire  cache_v__T_224_en; // @[icache.scala 91:18]
  wire  cache_v__T_225_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_225_addr; // @[icache.scala 91:18]
  wire  cache_v__T_225_mask; // @[icache.scala 91:18]
  wire  cache_v__T_225_en; // @[icache.scala 91:18]
  wire  cache_v__T_226_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_226_addr; // @[icache.scala 91:18]
  wire  cache_v__T_226_mask; // @[icache.scala 91:18]
  wire  cache_v__T_226_en; // @[icache.scala 91:18]
  wire  cache_v__T_227_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_227_addr; // @[icache.scala 91:18]
  wire  cache_v__T_227_mask; // @[icache.scala 91:18]
  wire  cache_v__T_227_en; // @[icache.scala 91:18]
  wire  cache_v__T_228_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_228_addr; // @[icache.scala 91:18]
  wire  cache_v__T_228_mask; // @[icache.scala 91:18]
  wire  cache_v__T_228_en; // @[icache.scala 91:18]
  wire  cache_v__T_229_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_229_addr; // @[icache.scala 91:18]
  wire  cache_v__T_229_mask; // @[icache.scala 91:18]
  wire  cache_v__T_229_en; // @[icache.scala 91:18]
  wire  cache_v__T_230_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_230_addr; // @[icache.scala 91:18]
  wire  cache_v__T_230_mask; // @[icache.scala 91:18]
  wire  cache_v__T_230_en; // @[icache.scala 91:18]
  wire  cache_v__T_231_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_231_addr; // @[icache.scala 91:18]
  wire  cache_v__T_231_mask; // @[icache.scala 91:18]
  wire  cache_v__T_231_en; // @[icache.scala 91:18]
  wire  cache_v__T_232_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_232_addr; // @[icache.scala 91:18]
  wire  cache_v__T_232_mask; // @[icache.scala 91:18]
  wire  cache_v__T_232_en; // @[icache.scala 91:18]
  wire  cache_v__T_233_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_233_addr; // @[icache.scala 91:18]
  wire  cache_v__T_233_mask; // @[icache.scala 91:18]
  wire  cache_v__T_233_en; // @[icache.scala 91:18]
  wire  cache_v__T_234_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_234_addr; // @[icache.scala 91:18]
  wire  cache_v__T_234_mask; // @[icache.scala 91:18]
  wire  cache_v__T_234_en; // @[icache.scala 91:18]
  wire  cache_v__T_235_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_235_addr; // @[icache.scala 91:18]
  wire  cache_v__T_235_mask; // @[icache.scala 91:18]
  wire  cache_v__T_235_en; // @[icache.scala 91:18]
  wire  cache_v__T_236_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_236_addr; // @[icache.scala 91:18]
  wire  cache_v__T_236_mask; // @[icache.scala 91:18]
  wire  cache_v__T_236_en; // @[icache.scala 91:18]
  wire  cache_v__T_237_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_237_addr; // @[icache.scala 91:18]
  wire  cache_v__T_237_mask; // @[icache.scala 91:18]
  wire  cache_v__T_237_en; // @[icache.scala 91:18]
  wire  cache_v__T_238_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_238_addr; // @[icache.scala 91:18]
  wire  cache_v__T_238_mask; // @[icache.scala 91:18]
  wire  cache_v__T_238_en; // @[icache.scala 91:18]
  wire  cache_v__T_239_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_239_addr; // @[icache.scala 91:18]
  wire  cache_v__T_239_mask; // @[icache.scala 91:18]
  wire  cache_v__T_239_en; // @[icache.scala 91:18]
  wire  cache_v__T_240_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_240_addr; // @[icache.scala 91:18]
  wire  cache_v__T_240_mask; // @[icache.scala 91:18]
  wire  cache_v__T_240_en; // @[icache.scala 91:18]
  wire  cache_v__T_241_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_241_addr; // @[icache.scala 91:18]
  wire  cache_v__T_241_mask; // @[icache.scala 91:18]
  wire  cache_v__T_241_en; // @[icache.scala 91:18]
  wire  cache_v__T_242_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_242_addr; // @[icache.scala 91:18]
  wire  cache_v__T_242_mask; // @[icache.scala 91:18]
  wire  cache_v__T_242_en; // @[icache.scala 91:18]
  wire  cache_v__T_243_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_243_addr; // @[icache.scala 91:18]
  wire  cache_v__T_243_mask; // @[icache.scala 91:18]
  wire  cache_v__T_243_en; // @[icache.scala 91:18]
  wire  cache_v__T_244_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_244_addr; // @[icache.scala 91:18]
  wire  cache_v__T_244_mask; // @[icache.scala 91:18]
  wire  cache_v__T_244_en; // @[icache.scala 91:18]
  wire  cache_v__T_245_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_245_addr; // @[icache.scala 91:18]
  wire  cache_v__T_245_mask; // @[icache.scala 91:18]
  wire  cache_v__T_245_en; // @[icache.scala 91:18]
  wire  cache_v__T_246_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_246_addr; // @[icache.scala 91:18]
  wire  cache_v__T_246_mask; // @[icache.scala 91:18]
  wire  cache_v__T_246_en; // @[icache.scala 91:18]
  wire  cache_v__T_247_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_247_addr; // @[icache.scala 91:18]
  wire  cache_v__T_247_mask; // @[icache.scala 91:18]
  wire  cache_v__T_247_en; // @[icache.scala 91:18]
  wire  cache_v__T_248_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_248_addr; // @[icache.scala 91:18]
  wire  cache_v__T_248_mask; // @[icache.scala 91:18]
  wire  cache_v__T_248_en; // @[icache.scala 91:18]
  wire  cache_v__T_249_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_249_addr; // @[icache.scala 91:18]
  wire  cache_v__T_249_mask; // @[icache.scala 91:18]
  wire  cache_v__T_249_en; // @[icache.scala 91:18]
  wire  cache_v__T_250_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_250_addr; // @[icache.scala 91:18]
  wire  cache_v__T_250_mask; // @[icache.scala 91:18]
  wire  cache_v__T_250_en; // @[icache.scala 91:18]
  wire  cache_v__T_251_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_251_addr; // @[icache.scala 91:18]
  wire  cache_v__T_251_mask; // @[icache.scala 91:18]
  wire  cache_v__T_251_en; // @[icache.scala 91:18]
  wire  cache_v__T_252_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_252_addr; // @[icache.scala 91:18]
  wire  cache_v__T_252_mask; // @[icache.scala 91:18]
  wire  cache_v__T_252_en; // @[icache.scala 91:18]
  wire  cache_v__T_253_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_253_addr; // @[icache.scala 91:18]
  wire  cache_v__T_253_mask; // @[icache.scala 91:18]
  wire  cache_v__T_253_en; // @[icache.scala 91:18]
  wire  cache_v__T_254_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_254_addr; // @[icache.scala 91:18]
  wire  cache_v__T_254_mask; // @[icache.scala 91:18]
  wire  cache_v__T_254_en; // @[icache.scala 91:18]
  wire  cache_v__T_255_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_255_addr; // @[icache.scala 91:18]
  wire  cache_v__T_255_mask; // @[icache.scala 91:18]
  wire  cache_v__T_255_en; // @[icache.scala 91:18]
  wire  cache_v__T_256_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_256_addr; // @[icache.scala 91:18]
  wire  cache_v__T_256_mask; // @[icache.scala 91:18]
  wire  cache_v__T_256_en; // @[icache.scala 91:18]
  wire  cache_v__T_257_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_257_addr; // @[icache.scala 91:18]
  wire  cache_v__T_257_mask; // @[icache.scala 91:18]
  wire  cache_v__T_257_en; // @[icache.scala 91:18]
  wire  cache_v__T_258_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_258_addr; // @[icache.scala 91:18]
  wire  cache_v__T_258_mask; // @[icache.scala 91:18]
  wire  cache_v__T_258_en; // @[icache.scala 91:18]
  wire  cache_v__T_259_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_259_addr; // @[icache.scala 91:18]
  wire  cache_v__T_259_mask; // @[icache.scala 91:18]
  wire  cache_v__T_259_en; // @[icache.scala 91:18]
  wire  cache_v__T_260_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_260_addr; // @[icache.scala 91:18]
  wire  cache_v__T_260_mask; // @[icache.scala 91:18]
  wire  cache_v__T_260_en; // @[icache.scala 91:18]
  wire  cache_v__T_261_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_261_addr; // @[icache.scala 91:18]
  wire  cache_v__T_261_mask; // @[icache.scala 91:18]
  wire  cache_v__T_261_en; // @[icache.scala 91:18]
  wire  cache_v__T_262_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_262_addr; // @[icache.scala 91:18]
  wire  cache_v__T_262_mask; // @[icache.scala 91:18]
  wire  cache_v__T_262_en; // @[icache.scala 91:18]
  wire  cache_v__T_263_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_263_addr; // @[icache.scala 91:18]
  wire  cache_v__T_263_mask; // @[icache.scala 91:18]
  wire  cache_v__T_263_en; // @[icache.scala 91:18]
  wire  cache_v__T_264_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_264_addr; // @[icache.scala 91:18]
  wire  cache_v__T_264_mask; // @[icache.scala 91:18]
  wire  cache_v__T_264_en; // @[icache.scala 91:18]
  wire  cache_v__T_265_data; // @[icache.scala 91:18]
  wire [7:0] cache_v__T_265_addr; // @[icache.scala 91:18]
  wire  cache_v__T_265_mask; // @[icache.scala 91:18]
  wire  cache_v__T_265_en; // @[icache.scala 91:18]
  wire  cache_v_s1_entry_w_data; // @[icache.scala 91:18]
  wire [7:0] cache_v_s1_entry_w_addr; // @[icache.scala 91:18]
  wire  cache_v_s1_entry_w_mask; // @[icache.scala 91:18]
  wire  cache_v_s1_entry_w_en; // @[icache.scala 91:18]
  reg [23:0] cache_tag [0:255]; // @[icache.scala 91:18]
  reg [31:0] _RAND_1;
  wire [23:0] cache_tag_s1_entry_r_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag_s1_entry_r_addr; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_8_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_8_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_8_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_8_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_10_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_10_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_10_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_10_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_11_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_11_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_11_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_11_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_12_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_12_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_12_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_12_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_13_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_13_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_13_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_13_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_14_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_14_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_14_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_14_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_15_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_15_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_15_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_15_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_16_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_16_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_16_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_16_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_17_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_17_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_17_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_17_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_18_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_18_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_18_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_18_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_19_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_19_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_19_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_19_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_20_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_20_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_20_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_20_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_21_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_21_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_21_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_21_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_22_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_22_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_22_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_22_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_23_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_23_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_23_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_23_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_24_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_24_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_24_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_24_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_25_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_25_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_25_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_25_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_26_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_26_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_26_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_26_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_27_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_27_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_27_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_27_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_28_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_28_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_28_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_28_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_29_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_29_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_29_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_29_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_30_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_30_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_30_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_30_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_31_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_31_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_31_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_31_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_32_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_32_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_32_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_32_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_33_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_33_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_33_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_33_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_34_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_34_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_34_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_34_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_35_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_35_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_35_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_35_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_36_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_36_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_36_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_36_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_37_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_37_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_37_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_37_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_38_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_38_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_38_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_38_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_39_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_39_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_39_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_39_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_40_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_40_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_40_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_40_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_41_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_41_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_41_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_41_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_42_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_42_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_42_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_42_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_43_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_43_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_43_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_43_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_44_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_44_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_44_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_44_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_45_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_45_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_45_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_45_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_46_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_46_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_46_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_46_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_47_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_47_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_47_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_47_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_48_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_48_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_48_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_48_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_49_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_49_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_49_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_49_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_50_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_50_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_50_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_50_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_51_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_51_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_51_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_51_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_52_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_52_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_52_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_52_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_53_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_53_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_53_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_53_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_54_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_54_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_54_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_54_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_55_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_55_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_55_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_55_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_56_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_56_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_56_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_56_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_57_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_57_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_57_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_57_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_58_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_58_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_58_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_58_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_59_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_59_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_59_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_59_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_60_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_60_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_60_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_60_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_61_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_61_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_61_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_61_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_62_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_62_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_62_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_62_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_63_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_63_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_63_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_63_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_64_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_64_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_64_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_64_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_65_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_65_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_65_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_65_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_66_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_66_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_66_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_66_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_67_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_67_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_67_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_67_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_68_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_68_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_68_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_68_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_69_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_69_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_69_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_69_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_70_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_70_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_70_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_70_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_71_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_71_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_71_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_71_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_72_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_72_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_72_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_72_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_73_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_73_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_73_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_73_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_74_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_74_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_74_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_74_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_75_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_75_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_75_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_75_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_76_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_76_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_76_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_76_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_77_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_77_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_77_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_77_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_78_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_78_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_78_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_78_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_79_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_79_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_79_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_79_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_80_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_80_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_80_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_80_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_81_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_81_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_81_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_81_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_82_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_82_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_82_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_82_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_83_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_83_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_83_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_83_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_84_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_84_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_84_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_84_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_85_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_85_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_85_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_85_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_86_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_86_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_86_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_86_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_87_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_87_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_87_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_87_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_88_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_88_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_88_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_88_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_89_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_89_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_89_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_89_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_90_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_90_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_90_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_90_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_91_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_91_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_91_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_91_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_92_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_92_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_92_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_92_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_93_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_93_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_93_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_93_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_94_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_94_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_94_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_94_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_95_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_95_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_95_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_95_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_96_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_96_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_96_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_96_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_97_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_97_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_97_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_97_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_98_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_98_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_98_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_98_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_99_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_99_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_99_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_99_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_100_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_100_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_100_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_100_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_101_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_101_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_101_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_101_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_102_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_102_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_102_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_102_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_103_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_103_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_103_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_103_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_104_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_104_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_104_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_104_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_105_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_105_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_105_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_105_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_106_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_106_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_106_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_106_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_107_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_107_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_107_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_107_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_108_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_108_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_108_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_108_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_109_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_109_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_109_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_109_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_110_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_110_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_110_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_110_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_111_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_111_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_111_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_111_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_112_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_112_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_112_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_112_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_113_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_113_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_113_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_113_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_114_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_114_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_114_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_114_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_115_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_115_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_115_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_115_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_116_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_116_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_116_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_116_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_117_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_117_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_117_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_117_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_118_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_118_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_118_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_118_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_119_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_119_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_119_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_119_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_120_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_120_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_120_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_120_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_121_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_121_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_121_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_121_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_122_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_122_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_122_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_122_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_123_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_123_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_123_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_123_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_124_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_124_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_124_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_124_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_125_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_125_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_125_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_125_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_126_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_126_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_126_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_126_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_127_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_127_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_127_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_127_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_128_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_128_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_128_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_128_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_129_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_129_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_129_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_129_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_130_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_130_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_130_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_130_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_131_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_131_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_131_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_131_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_132_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_132_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_132_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_132_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_133_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_133_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_133_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_133_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_134_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_134_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_134_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_134_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_135_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_135_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_135_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_135_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_136_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_136_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_136_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_136_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_137_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_137_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_137_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_137_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_138_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_138_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_138_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_138_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_139_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_139_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_139_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_139_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_140_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_140_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_140_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_140_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_141_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_141_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_141_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_141_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_142_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_142_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_142_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_142_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_143_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_143_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_143_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_143_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_144_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_144_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_144_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_144_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_145_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_145_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_145_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_145_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_146_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_146_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_146_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_146_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_147_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_147_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_147_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_147_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_148_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_148_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_148_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_148_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_149_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_149_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_149_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_149_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_150_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_150_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_150_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_150_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_151_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_151_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_151_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_151_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_152_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_152_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_152_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_152_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_153_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_153_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_153_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_153_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_154_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_154_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_154_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_154_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_155_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_155_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_155_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_155_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_156_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_156_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_156_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_156_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_157_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_157_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_157_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_157_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_158_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_158_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_158_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_158_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_159_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_159_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_159_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_159_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_160_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_160_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_160_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_160_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_161_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_161_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_161_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_161_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_162_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_162_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_162_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_162_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_163_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_163_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_163_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_163_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_164_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_164_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_164_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_164_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_165_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_165_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_165_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_165_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_166_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_166_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_166_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_166_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_167_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_167_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_167_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_167_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_168_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_168_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_168_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_168_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_169_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_169_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_169_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_169_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_170_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_170_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_170_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_170_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_171_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_171_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_171_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_171_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_172_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_172_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_172_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_172_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_173_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_173_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_173_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_173_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_174_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_174_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_174_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_174_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_175_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_175_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_175_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_175_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_176_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_176_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_176_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_176_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_177_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_177_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_177_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_177_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_178_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_178_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_178_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_178_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_179_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_179_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_179_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_179_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_180_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_180_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_180_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_180_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_181_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_181_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_181_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_181_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_182_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_182_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_182_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_182_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_183_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_183_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_183_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_183_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_184_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_184_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_184_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_184_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_185_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_185_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_185_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_185_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_186_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_186_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_186_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_186_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_187_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_187_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_187_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_187_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_188_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_188_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_188_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_188_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_189_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_189_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_189_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_189_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_190_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_190_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_190_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_190_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_191_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_191_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_191_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_191_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_192_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_192_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_192_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_192_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_193_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_193_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_193_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_193_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_194_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_194_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_194_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_194_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_195_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_195_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_195_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_195_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_196_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_196_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_196_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_196_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_197_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_197_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_197_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_197_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_198_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_198_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_198_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_198_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_199_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_199_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_199_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_199_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_200_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_200_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_200_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_200_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_201_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_201_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_201_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_201_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_202_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_202_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_202_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_202_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_203_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_203_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_203_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_203_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_204_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_204_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_204_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_204_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_205_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_205_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_205_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_205_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_206_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_206_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_206_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_206_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_207_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_207_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_207_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_207_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_208_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_208_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_208_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_208_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_209_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_209_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_209_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_209_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_210_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_210_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_210_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_210_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_211_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_211_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_211_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_211_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_212_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_212_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_212_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_212_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_213_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_213_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_213_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_213_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_214_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_214_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_214_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_214_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_215_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_215_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_215_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_215_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_216_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_216_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_216_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_216_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_217_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_217_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_217_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_217_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_218_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_218_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_218_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_218_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_219_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_219_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_219_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_219_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_220_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_220_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_220_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_220_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_221_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_221_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_221_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_221_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_222_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_222_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_222_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_222_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_223_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_223_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_223_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_223_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_224_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_224_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_224_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_224_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_225_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_225_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_225_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_225_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_226_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_226_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_226_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_226_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_227_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_227_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_227_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_227_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_228_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_228_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_228_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_228_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_229_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_229_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_229_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_229_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_230_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_230_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_230_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_230_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_231_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_231_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_231_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_231_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_232_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_232_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_232_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_232_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_233_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_233_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_233_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_233_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_234_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_234_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_234_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_234_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_235_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_235_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_235_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_235_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_236_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_236_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_236_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_236_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_237_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_237_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_237_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_237_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_238_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_238_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_238_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_238_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_239_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_239_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_239_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_239_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_240_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_240_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_240_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_240_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_241_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_241_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_241_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_241_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_242_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_242_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_242_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_242_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_243_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_243_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_243_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_243_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_244_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_244_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_244_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_244_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_245_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_245_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_245_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_245_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_246_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_246_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_246_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_246_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_247_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_247_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_247_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_247_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_248_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_248_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_248_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_248_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_249_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_249_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_249_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_249_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_250_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_250_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_250_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_250_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_251_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_251_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_251_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_251_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_252_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_252_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_252_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_252_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_253_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_253_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_253_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_253_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_254_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_254_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_254_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_254_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_255_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_255_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_255_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_255_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_256_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_256_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_256_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_256_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_257_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_257_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_257_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_257_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_258_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_258_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_258_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_258_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_259_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_259_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_259_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_259_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_260_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_260_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_260_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_260_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_261_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_261_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_261_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_261_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_262_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_262_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_262_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_262_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_263_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_263_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_263_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_263_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_264_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_264_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_264_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_264_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag__T_265_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag__T_265_addr; // @[icache.scala 91:18]
  wire  cache_tag__T_265_mask; // @[icache.scala 91:18]
  wire  cache_tag__T_265_en; // @[icache.scala 91:18]
  wire [23:0] cache_tag_s1_entry_w_data; // @[icache.scala 91:18]
  wire [7:0] cache_tag_s1_entry_w_addr; // @[icache.scala 91:18]
  wire  cache_tag_s1_entry_w_mask; // @[icache.scala 91:18]
  wire  cache_tag_s1_entry_w_en; // @[icache.scala 91:18]
  reg [31:0] cache_data [0:255]; // @[icache.scala 91:18]
  reg [31:0] _RAND_2;
  wire [31:0] cache_data_s1_entry_r_data; // @[icache.scala 91:18]
  wire [7:0] cache_data_s1_entry_r_addr; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_8_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_8_addr; // @[icache.scala 91:18]
  wire  cache_data__T_8_mask; // @[icache.scala 91:18]
  wire  cache_data__T_8_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_10_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_10_addr; // @[icache.scala 91:18]
  wire  cache_data__T_10_mask; // @[icache.scala 91:18]
  wire  cache_data__T_10_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_11_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_11_addr; // @[icache.scala 91:18]
  wire  cache_data__T_11_mask; // @[icache.scala 91:18]
  wire  cache_data__T_11_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_12_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_12_addr; // @[icache.scala 91:18]
  wire  cache_data__T_12_mask; // @[icache.scala 91:18]
  wire  cache_data__T_12_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_13_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_13_addr; // @[icache.scala 91:18]
  wire  cache_data__T_13_mask; // @[icache.scala 91:18]
  wire  cache_data__T_13_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_14_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_14_addr; // @[icache.scala 91:18]
  wire  cache_data__T_14_mask; // @[icache.scala 91:18]
  wire  cache_data__T_14_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_15_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_15_addr; // @[icache.scala 91:18]
  wire  cache_data__T_15_mask; // @[icache.scala 91:18]
  wire  cache_data__T_15_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_16_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_16_addr; // @[icache.scala 91:18]
  wire  cache_data__T_16_mask; // @[icache.scala 91:18]
  wire  cache_data__T_16_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_17_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_17_addr; // @[icache.scala 91:18]
  wire  cache_data__T_17_mask; // @[icache.scala 91:18]
  wire  cache_data__T_17_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_18_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_18_addr; // @[icache.scala 91:18]
  wire  cache_data__T_18_mask; // @[icache.scala 91:18]
  wire  cache_data__T_18_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_19_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_19_addr; // @[icache.scala 91:18]
  wire  cache_data__T_19_mask; // @[icache.scala 91:18]
  wire  cache_data__T_19_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_20_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_20_addr; // @[icache.scala 91:18]
  wire  cache_data__T_20_mask; // @[icache.scala 91:18]
  wire  cache_data__T_20_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_21_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_21_addr; // @[icache.scala 91:18]
  wire  cache_data__T_21_mask; // @[icache.scala 91:18]
  wire  cache_data__T_21_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_22_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_22_addr; // @[icache.scala 91:18]
  wire  cache_data__T_22_mask; // @[icache.scala 91:18]
  wire  cache_data__T_22_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_23_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_23_addr; // @[icache.scala 91:18]
  wire  cache_data__T_23_mask; // @[icache.scala 91:18]
  wire  cache_data__T_23_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_24_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_24_addr; // @[icache.scala 91:18]
  wire  cache_data__T_24_mask; // @[icache.scala 91:18]
  wire  cache_data__T_24_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_25_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_25_addr; // @[icache.scala 91:18]
  wire  cache_data__T_25_mask; // @[icache.scala 91:18]
  wire  cache_data__T_25_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_26_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_26_addr; // @[icache.scala 91:18]
  wire  cache_data__T_26_mask; // @[icache.scala 91:18]
  wire  cache_data__T_26_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_27_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_27_addr; // @[icache.scala 91:18]
  wire  cache_data__T_27_mask; // @[icache.scala 91:18]
  wire  cache_data__T_27_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_28_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_28_addr; // @[icache.scala 91:18]
  wire  cache_data__T_28_mask; // @[icache.scala 91:18]
  wire  cache_data__T_28_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_29_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_29_addr; // @[icache.scala 91:18]
  wire  cache_data__T_29_mask; // @[icache.scala 91:18]
  wire  cache_data__T_29_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_30_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_30_addr; // @[icache.scala 91:18]
  wire  cache_data__T_30_mask; // @[icache.scala 91:18]
  wire  cache_data__T_30_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_31_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_31_addr; // @[icache.scala 91:18]
  wire  cache_data__T_31_mask; // @[icache.scala 91:18]
  wire  cache_data__T_31_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_32_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_32_addr; // @[icache.scala 91:18]
  wire  cache_data__T_32_mask; // @[icache.scala 91:18]
  wire  cache_data__T_32_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_33_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_33_addr; // @[icache.scala 91:18]
  wire  cache_data__T_33_mask; // @[icache.scala 91:18]
  wire  cache_data__T_33_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_34_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_34_addr; // @[icache.scala 91:18]
  wire  cache_data__T_34_mask; // @[icache.scala 91:18]
  wire  cache_data__T_34_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_35_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_35_addr; // @[icache.scala 91:18]
  wire  cache_data__T_35_mask; // @[icache.scala 91:18]
  wire  cache_data__T_35_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_36_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_36_addr; // @[icache.scala 91:18]
  wire  cache_data__T_36_mask; // @[icache.scala 91:18]
  wire  cache_data__T_36_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_37_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_37_addr; // @[icache.scala 91:18]
  wire  cache_data__T_37_mask; // @[icache.scala 91:18]
  wire  cache_data__T_37_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_38_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_38_addr; // @[icache.scala 91:18]
  wire  cache_data__T_38_mask; // @[icache.scala 91:18]
  wire  cache_data__T_38_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_39_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_39_addr; // @[icache.scala 91:18]
  wire  cache_data__T_39_mask; // @[icache.scala 91:18]
  wire  cache_data__T_39_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_40_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_40_addr; // @[icache.scala 91:18]
  wire  cache_data__T_40_mask; // @[icache.scala 91:18]
  wire  cache_data__T_40_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_41_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_41_addr; // @[icache.scala 91:18]
  wire  cache_data__T_41_mask; // @[icache.scala 91:18]
  wire  cache_data__T_41_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_42_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_42_addr; // @[icache.scala 91:18]
  wire  cache_data__T_42_mask; // @[icache.scala 91:18]
  wire  cache_data__T_42_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_43_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_43_addr; // @[icache.scala 91:18]
  wire  cache_data__T_43_mask; // @[icache.scala 91:18]
  wire  cache_data__T_43_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_44_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_44_addr; // @[icache.scala 91:18]
  wire  cache_data__T_44_mask; // @[icache.scala 91:18]
  wire  cache_data__T_44_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_45_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_45_addr; // @[icache.scala 91:18]
  wire  cache_data__T_45_mask; // @[icache.scala 91:18]
  wire  cache_data__T_45_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_46_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_46_addr; // @[icache.scala 91:18]
  wire  cache_data__T_46_mask; // @[icache.scala 91:18]
  wire  cache_data__T_46_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_47_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_47_addr; // @[icache.scala 91:18]
  wire  cache_data__T_47_mask; // @[icache.scala 91:18]
  wire  cache_data__T_47_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_48_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_48_addr; // @[icache.scala 91:18]
  wire  cache_data__T_48_mask; // @[icache.scala 91:18]
  wire  cache_data__T_48_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_49_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_49_addr; // @[icache.scala 91:18]
  wire  cache_data__T_49_mask; // @[icache.scala 91:18]
  wire  cache_data__T_49_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_50_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_50_addr; // @[icache.scala 91:18]
  wire  cache_data__T_50_mask; // @[icache.scala 91:18]
  wire  cache_data__T_50_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_51_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_51_addr; // @[icache.scala 91:18]
  wire  cache_data__T_51_mask; // @[icache.scala 91:18]
  wire  cache_data__T_51_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_52_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_52_addr; // @[icache.scala 91:18]
  wire  cache_data__T_52_mask; // @[icache.scala 91:18]
  wire  cache_data__T_52_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_53_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_53_addr; // @[icache.scala 91:18]
  wire  cache_data__T_53_mask; // @[icache.scala 91:18]
  wire  cache_data__T_53_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_54_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_54_addr; // @[icache.scala 91:18]
  wire  cache_data__T_54_mask; // @[icache.scala 91:18]
  wire  cache_data__T_54_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_55_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_55_addr; // @[icache.scala 91:18]
  wire  cache_data__T_55_mask; // @[icache.scala 91:18]
  wire  cache_data__T_55_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_56_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_56_addr; // @[icache.scala 91:18]
  wire  cache_data__T_56_mask; // @[icache.scala 91:18]
  wire  cache_data__T_56_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_57_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_57_addr; // @[icache.scala 91:18]
  wire  cache_data__T_57_mask; // @[icache.scala 91:18]
  wire  cache_data__T_57_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_58_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_58_addr; // @[icache.scala 91:18]
  wire  cache_data__T_58_mask; // @[icache.scala 91:18]
  wire  cache_data__T_58_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_59_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_59_addr; // @[icache.scala 91:18]
  wire  cache_data__T_59_mask; // @[icache.scala 91:18]
  wire  cache_data__T_59_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_60_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_60_addr; // @[icache.scala 91:18]
  wire  cache_data__T_60_mask; // @[icache.scala 91:18]
  wire  cache_data__T_60_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_61_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_61_addr; // @[icache.scala 91:18]
  wire  cache_data__T_61_mask; // @[icache.scala 91:18]
  wire  cache_data__T_61_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_62_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_62_addr; // @[icache.scala 91:18]
  wire  cache_data__T_62_mask; // @[icache.scala 91:18]
  wire  cache_data__T_62_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_63_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_63_addr; // @[icache.scala 91:18]
  wire  cache_data__T_63_mask; // @[icache.scala 91:18]
  wire  cache_data__T_63_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_64_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_64_addr; // @[icache.scala 91:18]
  wire  cache_data__T_64_mask; // @[icache.scala 91:18]
  wire  cache_data__T_64_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_65_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_65_addr; // @[icache.scala 91:18]
  wire  cache_data__T_65_mask; // @[icache.scala 91:18]
  wire  cache_data__T_65_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_66_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_66_addr; // @[icache.scala 91:18]
  wire  cache_data__T_66_mask; // @[icache.scala 91:18]
  wire  cache_data__T_66_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_67_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_67_addr; // @[icache.scala 91:18]
  wire  cache_data__T_67_mask; // @[icache.scala 91:18]
  wire  cache_data__T_67_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_68_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_68_addr; // @[icache.scala 91:18]
  wire  cache_data__T_68_mask; // @[icache.scala 91:18]
  wire  cache_data__T_68_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_69_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_69_addr; // @[icache.scala 91:18]
  wire  cache_data__T_69_mask; // @[icache.scala 91:18]
  wire  cache_data__T_69_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_70_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_70_addr; // @[icache.scala 91:18]
  wire  cache_data__T_70_mask; // @[icache.scala 91:18]
  wire  cache_data__T_70_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_71_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_71_addr; // @[icache.scala 91:18]
  wire  cache_data__T_71_mask; // @[icache.scala 91:18]
  wire  cache_data__T_71_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_72_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_72_addr; // @[icache.scala 91:18]
  wire  cache_data__T_72_mask; // @[icache.scala 91:18]
  wire  cache_data__T_72_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_73_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_73_addr; // @[icache.scala 91:18]
  wire  cache_data__T_73_mask; // @[icache.scala 91:18]
  wire  cache_data__T_73_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_74_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_74_addr; // @[icache.scala 91:18]
  wire  cache_data__T_74_mask; // @[icache.scala 91:18]
  wire  cache_data__T_74_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_75_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_75_addr; // @[icache.scala 91:18]
  wire  cache_data__T_75_mask; // @[icache.scala 91:18]
  wire  cache_data__T_75_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_76_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_76_addr; // @[icache.scala 91:18]
  wire  cache_data__T_76_mask; // @[icache.scala 91:18]
  wire  cache_data__T_76_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_77_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_77_addr; // @[icache.scala 91:18]
  wire  cache_data__T_77_mask; // @[icache.scala 91:18]
  wire  cache_data__T_77_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_78_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_78_addr; // @[icache.scala 91:18]
  wire  cache_data__T_78_mask; // @[icache.scala 91:18]
  wire  cache_data__T_78_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_79_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_79_addr; // @[icache.scala 91:18]
  wire  cache_data__T_79_mask; // @[icache.scala 91:18]
  wire  cache_data__T_79_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_80_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_80_addr; // @[icache.scala 91:18]
  wire  cache_data__T_80_mask; // @[icache.scala 91:18]
  wire  cache_data__T_80_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_81_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_81_addr; // @[icache.scala 91:18]
  wire  cache_data__T_81_mask; // @[icache.scala 91:18]
  wire  cache_data__T_81_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_82_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_82_addr; // @[icache.scala 91:18]
  wire  cache_data__T_82_mask; // @[icache.scala 91:18]
  wire  cache_data__T_82_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_83_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_83_addr; // @[icache.scala 91:18]
  wire  cache_data__T_83_mask; // @[icache.scala 91:18]
  wire  cache_data__T_83_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_84_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_84_addr; // @[icache.scala 91:18]
  wire  cache_data__T_84_mask; // @[icache.scala 91:18]
  wire  cache_data__T_84_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_85_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_85_addr; // @[icache.scala 91:18]
  wire  cache_data__T_85_mask; // @[icache.scala 91:18]
  wire  cache_data__T_85_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_86_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_86_addr; // @[icache.scala 91:18]
  wire  cache_data__T_86_mask; // @[icache.scala 91:18]
  wire  cache_data__T_86_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_87_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_87_addr; // @[icache.scala 91:18]
  wire  cache_data__T_87_mask; // @[icache.scala 91:18]
  wire  cache_data__T_87_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_88_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_88_addr; // @[icache.scala 91:18]
  wire  cache_data__T_88_mask; // @[icache.scala 91:18]
  wire  cache_data__T_88_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_89_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_89_addr; // @[icache.scala 91:18]
  wire  cache_data__T_89_mask; // @[icache.scala 91:18]
  wire  cache_data__T_89_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_90_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_90_addr; // @[icache.scala 91:18]
  wire  cache_data__T_90_mask; // @[icache.scala 91:18]
  wire  cache_data__T_90_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_91_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_91_addr; // @[icache.scala 91:18]
  wire  cache_data__T_91_mask; // @[icache.scala 91:18]
  wire  cache_data__T_91_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_92_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_92_addr; // @[icache.scala 91:18]
  wire  cache_data__T_92_mask; // @[icache.scala 91:18]
  wire  cache_data__T_92_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_93_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_93_addr; // @[icache.scala 91:18]
  wire  cache_data__T_93_mask; // @[icache.scala 91:18]
  wire  cache_data__T_93_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_94_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_94_addr; // @[icache.scala 91:18]
  wire  cache_data__T_94_mask; // @[icache.scala 91:18]
  wire  cache_data__T_94_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_95_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_95_addr; // @[icache.scala 91:18]
  wire  cache_data__T_95_mask; // @[icache.scala 91:18]
  wire  cache_data__T_95_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_96_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_96_addr; // @[icache.scala 91:18]
  wire  cache_data__T_96_mask; // @[icache.scala 91:18]
  wire  cache_data__T_96_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_97_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_97_addr; // @[icache.scala 91:18]
  wire  cache_data__T_97_mask; // @[icache.scala 91:18]
  wire  cache_data__T_97_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_98_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_98_addr; // @[icache.scala 91:18]
  wire  cache_data__T_98_mask; // @[icache.scala 91:18]
  wire  cache_data__T_98_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_99_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_99_addr; // @[icache.scala 91:18]
  wire  cache_data__T_99_mask; // @[icache.scala 91:18]
  wire  cache_data__T_99_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_100_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_100_addr; // @[icache.scala 91:18]
  wire  cache_data__T_100_mask; // @[icache.scala 91:18]
  wire  cache_data__T_100_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_101_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_101_addr; // @[icache.scala 91:18]
  wire  cache_data__T_101_mask; // @[icache.scala 91:18]
  wire  cache_data__T_101_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_102_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_102_addr; // @[icache.scala 91:18]
  wire  cache_data__T_102_mask; // @[icache.scala 91:18]
  wire  cache_data__T_102_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_103_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_103_addr; // @[icache.scala 91:18]
  wire  cache_data__T_103_mask; // @[icache.scala 91:18]
  wire  cache_data__T_103_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_104_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_104_addr; // @[icache.scala 91:18]
  wire  cache_data__T_104_mask; // @[icache.scala 91:18]
  wire  cache_data__T_104_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_105_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_105_addr; // @[icache.scala 91:18]
  wire  cache_data__T_105_mask; // @[icache.scala 91:18]
  wire  cache_data__T_105_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_106_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_106_addr; // @[icache.scala 91:18]
  wire  cache_data__T_106_mask; // @[icache.scala 91:18]
  wire  cache_data__T_106_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_107_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_107_addr; // @[icache.scala 91:18]
  wire  cache_data__T_107_mask; // @[icache.scala 91:18]
  wire  cache_data__T_107_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_108_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_108_addr; // @[icache.scala 91:18]
  wire  cache_data__T_108_mask; // @[icache.scala 91:18]
  wire  cache_data__T_108_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_109_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_109_addr; // @[icache.scala 91:18]
  wire  cache_data__T_109_mask; // @[icache.scala 91:18]
  wire  cache_data__T_109_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_110_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_110_addr; // @[icache.scala 91:18]
  wire  cache_data__T_110_mask; // @[icache.scala 91:18]
  wire  cache_data__T_110_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_111_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_111_addr; // @[icache.scala 91:18]
  wire  cache_data__T_111_mask; // @[icache.scala 91:18]
  wire  cache_data__T_111_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_112_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_112_addr; // @[icache.scala 91:18]
  wire  cache_data__T_112_mask; // @[icache.scala 91:18]
  wire  cache_data__T_112_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_113_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_113_addr; // @[icache.scala 91:18]
  wire  cache_data__T_113_mask; // @[icache.scala 91:18]
  wire  cache_data__T_113_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_114_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_114_addr; // @[icache.scala 91:18]
  wire  cache_data__T_114_mask; // @[icache.scala 91:18]
  wire  cache_data__T_114_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_115_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_115_addr; // @[icache.scala 91:18]
  wire  cache_data__T_115_mask; // @[icache.scala 91:18]
  wire  cache_data__T_115_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_116_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_116_addr; // @[icache.scala 91:18]
  wire  cache_data__T_116_mask; // @[icache.scala 91:18]
  wire  cache_data__T_116_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_117_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_117_addr; // @[icache.scala 91:18]
  wire  cache_data__T_117_mask; // @[icache.scala 91:18]
  wire  cache_data__T_117_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_118_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_118_addr; // @[icache.scala 91:18]
  wire  cache_data__T_118_mask; // @[icache.scala 91:18]
  wire  cache_data__T_118_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_119_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_119_addr; // @[icache.scala 91:18]
  wire  cache_data__T_119_mask; // @[icache.scala 91:18]
  wire  cache_data__T_119_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_120_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_120_addr; // @[icache.scala 91:18]
  wire  cache_data__T_120_mask; // @[icache.scala 91:18]
  wire  cache_data__T_120_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_121_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_121_addr; // @[icache.scala 91:18]
  wire  cache_data__T_121_mask; // @[icache.scala 91:18]
  wire  cache_data__T_121_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_122_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_122_addr; // @[icache.scala 91:18]
  wire  cache_data__T_122_mask; // @[icache.scala 91:18]
  wire  cache_data__T_122_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_123_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_123_addr; // @[icache.scala 91:18]
  wire  cache_data__T_123_mask; // @[icache.scala 91:18]
  wire  cache_data__T_123_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_124_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_124_addr; // @[icache.scala 91:18]
  wire  cache_data__T_124_mask; // @[icache.scala 91:18]
  wire  cache_data__T_124_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_125_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_125_addr; // @[icache.scala 91:18]
  wire  cache_data__T_125_mask; // @[icache.scala 91:18]
  wire  cache_data__T_125_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_126_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_126_addr; // @[icache.scala 91:18]
  wire  cache_data__T_126_mask; // @[icache.scala 91:18]
  wire  cache_data__T_126_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_127_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_127_addr; // @[icache.scala 91:18]
  wire  cache_data__T_127_mask; // @[icache.scala 91:18]
  wire  cache_data__T_127_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_128_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_128_addr; // @[icache.scala 91:18]
  wire  cache_data__T_128_mask; // @[icache.scala 91:18]
  wire  cache_data__T_128_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_129_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_129_addr; // @[icache.scala 91:18]
  wire  cache_data__T_129_mask; // @[icache.scala 91:18]
  wire  cache_data__T_129_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_130_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_130_addr; // @[icache.scala 91:18]
  wire  cache_data__T_130_mask; // @[icache.scala 91:18]
  wire  cache_data__T_130_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_131_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_131_addr; // @[icache.scala 91:18]
  wire  cache_data__T_131_mask; // @[icache.scala 91:18]
  wire  cache_data__T_131_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_132_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_132_addr; // @[icache.scala 91:18]
  wire  cache_data__T_132_mask; // @[icache.scala 91:18]
  wire  cache_data__T_132_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_133_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_133_addr; // @[icache.scala 91:18]
  wire  cache_data__T_133_mask; // @[icache.scala 91:18]
  wire  cache_data__T_133_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_134_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_134_addr; // @[icache.scala 91:18]
  wire  cache_data__T_134_mask; // @[icache.scala 91:18]
  wire  cache_data__T_134_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_135_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_135_addr; // @[icache.scala 91:18]
  wire  cache_data__T_135_mask; // @[icache.scala 91:18]
  wire  cache_data__T_135_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_136_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_136_addr; // @[icache.scala 91:18]
  wire  cache_data__T_136_mask; // @[icache.scala 91:18]
  wire  cache_data__T_136_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_137_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_137_addr; // @[icache.scala 91:18]
  wire  cache_data__T_137_mask; // @[icache.scala 91:18]
  wire  cache_data__T_137_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_138_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_138_addr; // @[icache.scala 91:18]
  wire  cache_data__T_138_mask; // @[icache.scala 91:18]
  wire  cache_data__T_138_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_139_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_139_addr; // @[icache.scala 91:18]
  wire  cache_data__T_139_mask; // @[icache.scala 91:18]
  wire  cache_data__T_139_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_140_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_140_addr; // @[icache.scala 91:18]
  wire  cache_data__T_140_mask; // @[icache.scala 91:18]
  wire  cache_data__T_140_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_141_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_141_addr; // @[icache.scala 91:18]
  wire  cache_data__T_141_mask; // @[icache.scala 91:18]
  wire  cache_data__T_141_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_142_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_142_addr; // @[icache.scala 91:18]
  wire  cache_data__T_142_mask; // @[icache.scala 91:18]
  wire  cache_data__T_142_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_143_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_143_addr; // @[icache.scala 91:18]
  wire  cache_data__T_143_mask; // @[icache.scala 91:18]
  wire  cache_data__T_143_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_144_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_144_addr; // @[icache.scala 91:18]
  wire  cache_data__T_144_mask; // @[icache.scala 91:18]
  wire  cache_data__T_144_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_145_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_145_addr; // @[icache.scala 91:18]
  wire  cache_data__T_145_mask; // @[icache.scala 91:18]
  wire  cache_data__T_145_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_146_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_146_addr; // @[icache.scala 91:18]
  wire  cache_data__T_146_mask; // @[icache.scala 91:18]
  wire  cache_data__T_146_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_147_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_147_addr; // @[icache.scala 91:18]
  wire  cache_data__T_147_mask; // @[icache.scala 91:18]
  wire  cache_data__T_147_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_148_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_148_addr; // @[icache.scala 91:18]
  wire  cache_data__T_148_mask; // @[icache.scala 91:18]
  wire  cache_data__T_148_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_149_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_149_addr; // @[icache.scala 91:18]
  wire  cache_data__T_149_mask; // @[icache.scala 91:18]
  wire  cache_data__T_149_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_150_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_150_addr; // @[icache.scala 91:18]
  wire  cache_data__T_150_mask; // @[icache.scala 91:18]
  wire  cache_data__T_150_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_151_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_151_addr; // @[icache.scala 91:18]
  wire  cache_data__T_151_mask; // @[icache.scala 91:18]
  wire  cache_data__T_151_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_152_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_152_addr; // @[icache.scala 91:18]
  wire  cache_data__T_152_mask; // @[icache.scala 91:18]
  wire  cache_data__T_152_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_153_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_153_addr; // @[icache.scala 91:18]
  wire  cache_data__T_153_mask; // @[icache.scala 91:18]
  wire  cache_data__T_153_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_154_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_154_addr; // @[icache.scala 91:18]
  wire  cache_data__T_154_mask; // @[icache.scala 91:18]
  wire  cache_data__T_154_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_155_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_155_addr; // @[icache.scala 91:18]
  wire  cache_data__T_155_mask; // @[icache.scala 91:18]
  wire  cache_data__T_155_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_156_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_156_addr; // @[icache.scala 91:18]
  wire  cache_data__T_156_mask; // @[icache.scala 91:18]
  wire  cache_data__T_156_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_157_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_157_addr; // @[icache.scala 91:18]
  wire  cache_data__T_157_mask; // @[icache.scala 91:18]
  wire  cache_data__T_157_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_158_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_158_addr; // @[icache.scala 91:18]
  wire  cache_data__T_158_mask; // @[icache.scala 91:18]
  wire  cache_data__T_158_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_159_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_159_addr; // @[icache.scala 91:18]
  wire  cache_data__T_159_mask; // @[icache.scala 91:18]
  wire  cache_data__T_159_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_160_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_160_addr; // @[icache.scala 91:18]
  wire  cache_data__T_160_mask; // @[icache.scala 91:18]
  wire  cache_data__T_160_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_161_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_161_addr; // @[icache.scala 91:18]
  wire  cache_data__T_161_mask; // @[icache.scala 91:18]
  wire  cache_data__T_161_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_162_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_162_addr; // @[icache.scala 91:18]
  wire  cache_data__T_162_mask; // @[icache.scala 91:18]
  wire  cache_data__T_162_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_163_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_163_addr; // @[icache.scala 91:18]
  wire  cache_data__T_163_mask; // @[icache.scala 91:18]
  wire  cache_data__T_163_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_164_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_164_addr; // @[icache.scala 91:18]
  wire  cache_data__T_164_mask; // @[icache.scala 91:18]
  wire  cache_data__T_164_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_165_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_165_addr; // @[icache.scala 91:18]
  wire  cache_data__T_165_mask; // @[icache.scala 91:18]
  wire  cache_data__T_165_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_166_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_166_addr; // @[icache.scala 91:18]
  wire  cache_data__T_166_mask; // @[icache.scala 91:18]
  wire  cache_data__T_166_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_167_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_167_addr; // @[icache.scala 91:18]
  wire  cache_data__T_167_mask; // @[icache.scala 91:18]
  wire  cache_data__T_167_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_168_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_168_addr; // @[icache.scala 91:18]
  wire  cache_data__T_168_mask; // @[icache.scala 91:18]
  wire  cache_data__T_168_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_169_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_169_addr; // @[icache.scala 91:18]
  wire  cache_data__T_169_mask; // @[icache.scala 91:18]
  wire  cache_data__T_169_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_170_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_170_addr; // @[icache.scala 91:18]
  wire  cache_data__T_170_mask; // @[icache.scala 91:18]
  wire  cache_data__T_170_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_171_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_171_addr; // @[icache.scala 91:18]
  wire  cache_data__T_171_mask; // @[icache.scala 91:18]
  wire  cache_data__T_171_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_172_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_172_addr; // @[icache.scala 91:18]
  wire  cache_data__T_172_mask; // @[icache.scala 91:18]
  wire  cache_data__T_172_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_173_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_173_addr; // @[icache.scala 91:18]
  wire  cache_data__T_173_mask; // @[icache.scala 91:18]
  wire  cache_data__T_173_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_174_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_174_addr; // @[icache.scala 91:18]
  wire  cache_data__T_174_mask; // @[icache.scala 91:18]
  wire  cache_data__T_174_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_175_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_175_addr; // @[icache.scala 91:18]
  wire  cache_data__T_175_mask; // @[icache.scala 91:18]
  wire  cache_data__T_175_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_176_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_176_addr; // @[icache.scala 91:18]
  wire  cache_data__T_176_mask; // @[icache.scala 91:18]
  wire  cache_data__T_176_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_177_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_177_addr; // @[icache.scala 91:18]
  wire  cache_data__T_177_mask; // @[icache.scala 91:18]
  wire  cache_data__T_177_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_178_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_178_addr; // @[icache.scala 91:18]
  wire  cache_data__T_178_mask; // @[icache.scala 91:18]
  wire  cache_data__T_178_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_179_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_179_addr; // @[icache.scala 91:18]
  wire  cache_data__T_179_mask; // @[icache.scala 91:18]
  wire  cache_data__T_179_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_180_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_180_addr; // @[icache.scala 91:18]
  wire  cache_data__T_180_mask; // @[icache.scala 91:18]
  wire  cache_data__T_180_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_181_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_181_addr; // @[icache.scala 91:18]
  wire  cache_data__T_181_mask; // @[icache.scala 91:18]
  wire  cache_data__T_181_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_182_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_182_addr; // @[icache.scala 91:18]
  wire  cache_data__T_182_mask; // @[icache.scala 91:18]
  wire  cache_data__T_182_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_183_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_183_addr; // @[icache.scala 91:18]
  wire  cache_data__T_183_mask; // @[icache.scala 91:18]
  wire  cache_data__T_183_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_184_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_184_addr; // @[icache.scala 91:18]
  wire  cache_data__T_184_mask; // @[icache.scala 91:18]
  wire  cache_data__T_184_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_185_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_185_addr; // @[icache.scala 91:18]
  wire  cache_data__T_185_mask; // @[icache.scala 91:18]
  wire  cache_data__T_185_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_186_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_186_addr; // @[icache.scala 91:18]
  wire  cache_data__T_186_mask; // @[icache.scala 91:18]
  wire  cache_data__T_186_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_187_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_187_addr; // @[icache.scala 91:18]
  wire  cache_data__T_187_mask; // @[icache.scala 91:18]
  wire  cache_data__T_187_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_188_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_188_addr; // @[icache.scala 91:18]
  wire  cache_data__T_188_mask; // @[icache.scala 91:18]
  wire  cache_data__T_188_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_189_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_189_addr; // @[icache.scala 91:18]
  wire  cache_data__T_189_mask; // @[icache.scala 91:18]
  wire  cache_data__T_189_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_190_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_190_addr; // @[icache.scala 91:18]
  wire  cache_data__T_190_mask; // @[icache.scala 91:18]
  wire  cache_data__T_190_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_191_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_191_addr; // @[icache.scala 91:18]
  wire  cache_data__T_191_mask; // @[icache.scala 91:18]
  wire  cache_data__T_191_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_192_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_192_addr; // @[icache.scala 91:18]
  wire  cache_data__T_192_mask; // @[icache.scala 91:18]
  wire  cache_data__T_192_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_193_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_193_addr; // @[icache.scala 91:18]
  wire  cache_data__T_193_mask; // @[icache.scala 91:18]
  wire  cache_data__T_193_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_194_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_194_addr; // @[icache.scala 91:18]
  wire  cache_data__T_194_mask; // @[icache.scala 91:18]
  wire  cache_data__T_194_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_195_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_195_addr; // @[icache.scala 91:18]
  wire  cache_data__T_195_mask; // @[icache.scala 91:18]
  wire  cache_data__T_195_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_196_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_196_addr; // @[icache.scala 91:18]
  wire  cache_data__T_196_mask; // @[icache.scala 91:18]
  wire  cache_data__T_196_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_197_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_197_addr; // @[icache.scala 91:18]
  wire  cache_data__T_197_mask; // @[icache.scala 91:18]
  wire  cache_data__T_197_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_198_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_198_addr; // @[icache.scala 91:18]
  wire  cache_data__T_198_mask; // @[icache.scala 91:18]
  wire  cache_data__T_198_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_199_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_199_addr; // @[icache.scala 91:18]
  wire  cache_data__T_199_mask; // @[icache.scala 91:18]
  wire  cache_data__T_199_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_200_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_200_addr; // @[icache.scala 91:18]
  wire  cache_data__T_200_mask; // @[icache.scala 91:18]
  wire  cache_data__T_200_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_201_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_201_addr; // @[icache.scala 91:18]
  wire  cache_data__T_201_mask; // @[icache.scala 91:18]
  wire  cache_data__T_201_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_202_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_202_addr; // @[icache.scala 91:18]
  wire  cache_data__T_202_mask; // @[icache.scala 91:18]
  wire  cache_data__T_202_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_203_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_203_addr; // @[icache.scala 91:18]
  wire  cache_data__T_203_mask; // @[icache.scala 91:18]
  wire  cache_data__T_203_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_204_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_204_addr; // @[icache.scala 91:18]
  wire  cache_data__T_204_mask; // @[icache.scala 91:18]
  wire  cache_data__T_204_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_205_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_205_addr; // @[icache.scala 91:18]
  wire  cache_data__T_205_mask; // @[icache.scala 91:18]
  wire  cache_data__T_205_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_206_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_206_addr; // @[icache.scala 91:18]
  wire  cache_data__T_206_mask; // @[icache.scala 91:18]
  wire  cache_data__T_206_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_207_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_207_addr; // @[icache.scala 91:18]
  wire  cache_data__T_207_mask; // @[icache.scala 91:18]
  wire  cache_data__T_207_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_208_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_208_addr; // @[icache.scala 91:18]
  wire  cache_data__T_208_mask; // @[icache.scala 91:18]
  wire  cache_data__T_208_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_209_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_209_addr; // @[icache.scala 91:18]
  wire  cache_data__T_209_mask; // @[icache.scala 91:18]
  wire  cache_data__T_209_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_210_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_210_addr; // @[icache.scala 91:18]
  wire  cache_data__T_210_mask; // @[icache.scala 91:18]
  wire  cache_data__T_210_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_211_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_211_addr; // @[icache.scala 91:18]
  wire  cache_data__T_211_mask; // @[icache.scala 91:18]
  wire  cache_data__T_211_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_212_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_212_addr; // @[icache.scala 91:18]
  wire  cache_data__T_212_mask; // @[icache.scala 91:18]
  wire  cache_data__T_212_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_213_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_213_addr; // @[icache.scala 91:18]
  wire  cache_data__T_213_mask; // @[icache.scala 91:18]
  wire  cache_data__T_213_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_214_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_214_addr; // @[icache.scala 91:18]
  wire  cache_data__T_214_mask; // @[icache.scala 91:18]
  wire  cache_data__T_214_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_215_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_215_addr; // @[icache.scala 91:18]
  wire  cache_data__T_215_mask; // @[icache.scala 91:18]
  wire  cache_data__T_215_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_216_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_216_addr; // @[icache.scala 91:18]
  wire  cache_data__T_216_mask; // @[icache.scala 91:18]
  wire  cache_data__T_216_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_217_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_217_addr; // @[icache.scala 91:18]
  wire  cache_data__T_217_mask; // @[icache.scala 91:18]
  wire  cache_data__T_217_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_218_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_218_addr; // @[icache.scala 91:18]
  wire  cache_data__T_218_mask; // @[icache.scala 91:18]
  wire  cache_data__T_218_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_219_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_219_addr; // @[icache.scala 91:18]
  wire  cache_data__T_219_mask; // @[icache.scala 91:18]
  wire  cache_data__T_219_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_220_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_220_addr; // @[icache.scala 91:18]
  wire  cache_data__T_220_mask; // @[icache.scala 91:18]
  wire  cache_data__T_220_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_221_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_221_addr; // @[icache.scala 91:18]
  wire  cache_data__T_221_mask; // @[icache.scala 91:18]
  wire  cache_data__T_221_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_222_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_222_addr; // @[icache.scala 91:18]
  wire  cache_data__T_222_mask; // @[icache.scala 91:18]
  wire  cache_data__T_222_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_223_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_223_addr; // @[icache.scala 91:18]
  wire  cache_data__T_223_mask; // @[icache.scala 91:18]
  wire  cache_data__T_223_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_224_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_224_addr; // @[icache.scala 91:18]
  wire  cache_data__T_224_mask; // @[icache.scala 91:18]
  wire  cache_data__T_224_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_225_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_225_addr; // @[icache.scala 91:18]
  wire  cache_data__T_225_mask; // @[icache.scala 91:18]
  wire  cache_data__T_225_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_226_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_226_addr; // @[icache.scala 91:18]
  wire  cache_data__T_226_mask; // @[icache.scala 91:18]
  wire  cache_data__T_226_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_227_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_227_addr; // @[icache.scala 91:18]
  wire  cache_data__T_227_mask; // @[icache.scala 91:18]
  wire  cache_data__T_227_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_228_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_228_addr; // @[icache.scala 91:18]
  wire  cache_data__T_228_mask; // @[icache.scala 91:18]
  wire  cache_data__T_228_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_229_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_229_addr; // @[icache.scala 91:18]
  wire  cache_data__T_229_mask; // @[icache.scala 91:18]
  wire  cache_data__T_229_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_230_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_230_addr; // @[icache.scala 91:18]
  wire  cache_data__T_230_mask; // @[icache.scala 91:18]
  wire  cache_data__T_230_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_231_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_231_addr; // @[icache.scala 91:18]
  wire  cache_data__T_231_mask; // @[icache.scala 91:18]
  wire  cache_data__T_231_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_232_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_232_addr; // @[icache.scala 91:18]
  wire  cache_data__T_232_mask; // @[icache.scala 91:18]
  wire  cache_data__T_232_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_233_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_233_addr; // @[icache.scala 91:18]
  wire  cache_data__T_233_mask; // @[icache.scala 91:18]
  wire  cache_data__T_233_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_234_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_234_addr; // @[icache.scala 91:18]
  wire  cache_data__T_234_mask; // @[icache.scala 91:18]
  wire  cache_data__T_234_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_235_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_235_addr; // @[icache.scala 91:18]
  wire  cache_data__T_235_mask; // @[icache.scala 91:18]
  wire  cache_data__T_235_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_236_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_236_addr; // @[icache.scala 91:18]
  wire  cache_data__T_236_mask; // @[icache.scala 91:18]
  wire  cache_data__T_236_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_237_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_237_addr; // @[icache.scala 91:18]
  wire  cache_data__T_237_mask; // @[icache.scala 91:18]
  wire  cache_data__T_237_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_238_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_238_addr; // @[icache.scala 91:18]
  wire  cache_data__T_238_mask; // @[icache.scala 91:18]
  wire  cache_data__T_238_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_239_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_239_addr; // @[icache.scala 91:18]
  wire  cache_data__T_239_mask; // @[icache.scala 91:18]
  wire  cache_data__T_239_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_240_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_240_addr; // @[icache.scala 91:18]
  wire  cache_data__T_240_mask; // @[icache.scala 91:18]
  wire  cache_data__T_240_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_241_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_241_addr; // @[icache.scala 91:18]
  wire  cache_data__T_241_mask; // @[icache.scala 91:18]
  wire  cache_data__T_241_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_242_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_242_addr; // @[icache.scala 91:18]
  wire  cache_data__T_242_mask; // @[icache.scala 91:18]
  wire  cache_data__T_242_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_243_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_243_addr; // @[icache.scala 91:18]
  wire  cache_data__T_243_mask; // @[icache.scala 91:18]
  wire  cache_data__T_243_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_244_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_244_addr; // @[icache.scala 91:18]
  wire  cache_data__T_244_mask; // @[icache.scala 91:18]
  wire  cache_data__T_244_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_245_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_245_addr; // @[icache.scala 91:18]
  wire  cache_data__T_245_mask; // @[icache.scala 91:18]
  wire  cache_data__T_245_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_246_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_246_addr; // @[icache.scala 91:18]
  wire  cache_data__T_246_mask; // @[icache.scala 91:18]
  wire  cache_data__T_246_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_247_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_247_addr; // @[icache.scala 91:18]
  wire  cache_data__T_247_mask; // @[icache.scala 91:18]
  wire  cache_data__T_247_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_248_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_248_addr; // @[icache.scala 91:18]
  wire  cache_data__T_248_mask; // @[icache.scala 91:18]
  wire  cache_data__T_248_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_249_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_249_addr; // @[icache.scala 91:18]
  wire  cache_data__T_249_mask; // @[icache.scala 91:18]
  wire  cache_data__T_249_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_250_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_250_addr; // @[icache.scala 91:18]
  wire  cache_data__T_250_mask; // @[icache.scala 91:18]
  wire  cache_data__T_250_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_251_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_251_addr; // @[icache.scala 91:18]
  wire  cache_data__T_251_mask; // @[icache.scala 91:18]
  wire  cache_data__T_251_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_252_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_252_addr; // @[icache.scala 91:18]
  wire  cache_data__T_252_mask; // @[icache.scala 91:18]
  wire  cache_data__T_252_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_253_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_253_addr; // @[icache.scala 91:18]
  wire  cache_data__T_253_mask; // @[icache.scala 91:18]
  wire  cache_data__T_253_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_254_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_254_addr; // @[icache.scala 91:18]
  wire  cache_data__T_254_mask; // @[icache.scala 91:18]
  wire  cache_data__T_254_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_255_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_255_addr; // @[icache.scala 91:18]
  wire  cache_data__T_255_mask; // @[icache.scala 91:18]
  wire  cache_data__T_255_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_256_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_256_addr; // @[icache.scala 91:18]
  wire  cache_data__T_256_mask; // @[icache.scala 91:18]
  wire  cache_data__T_256_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_257_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_257_addr; // @[icache.scala 91:18]
  wire  cache_data__T_257_mask; // @[icache.scala 91:18]
  wire  cache_data__T_257_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_258_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_258_addr; // @[icache.scala 91:18]
  wire  cache_data__T_258_mask; // @[icache.scala 91:18]
  wire  cache_data__T_258_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_259_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_259_addr; // @[icache.scala 91:18]
  wire  cache_data__T_259_mask; // @[icache.scala 91:18]
  wire  cache_data__T_259_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_260_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_260_addr; // @[icache.scala 91:18]
  wire  cache_data__T_260_mask; // @[icache.scala 91:18]
  wire  cache_data__T_260_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_261_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_261_addr; // @[icache.scala 91:18]
  wire  cache_data__T_261_mask; // @[icache.scala 91:18]
  wire  cache_data__T_261_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_262_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_262_addr; // @[icache.scala 91:18]
  wire  cache_data__T_262_mask; // @[icache.scala 91:18]
  wire  cache_data__T_262_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_263_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_263_addr; // @[icache.scala 91:18]
  wire  cache_data__T_263_mask; // @[icache.scala 91:18]
  wire  cache_data__T_263_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_264_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_264_addr; // @[icache.scala 91:18]
  wire  cache_data__T_264_mask; // @[icache.scala 91:18]
  wire  cache_data__T_264_en; // @[icache.scala 91:18]
  wire [31:0] cache_data__T_265_data; // @[icache.scala 91:18]
  wire [7:0] cache_data__T_265_addr; // @[icache.scala 91:18]
  wire  cache_data__T_265_mask; // @[icache.scala 91:18]
  wire  cache_data__T_265_en; // @[icache.scala 91:18]
  wire [31:0] cache_data_s1_entry_w_data; // @[icache.scala 91:18]
  wire [7:0] cache_data_s1_entry_w_addr; // @[icache.scala 91:18]
  wire  cache_data_s1_entry_w_mask; // @[icache.scala 91:18]
  wire  cache_data_s1_entry_w_en; // @[icache.scala 91:18]
  wire  _T = ~io_ex_flush; // @[icache.scala 93:29]
  wire  _T_1 = io_control_valid & _T; // @[icache.scala 93:26]
  wire  _T_3 = io_control_bits_op == 3'h0; // @[icache.scala 97:30]
  wire  _T_4 = io_control_bits_op == 3'h4; // @[icache.scala 98:26]
  wire  _T_5 = _T_3 | _T_4; // @[icache.scala 97:53]
  wire [8:0] _T_6 = {1'h0,io_control_bits_addr[7:0]}; // @[Cat.scala 29:58]
  wire  flush = io_br_flush | io_ex_flush; // @[icache.scala 111:27]
  reg  s0_valid; // @[icache.scala 113:25]
  reg [31:0] _RAND_3;
  wire  _T_266 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  s0_in_is_cached; // @[Reg.scala 27:20]
  reg [31:0] _RAND_4;
  reg [31:0] s0_in_addr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_5;
  reg [1:0] s0_in_len; // @[Reg.scala 27:20]
  reg [31:0] _RAND_6;
  reg [3:0] s0_in_strb; // @[Reg.scala 27:20]
  reg [31:0] _RAND_7;
  reg [31:0] s1_in_addr; // @[Reg.scala 27:20]
  reg [31:0] _RAND_8;
  wire [23:0] s1_tag = s1_in_addr[31:8]; // @[icache.scala 90:30]
  wire  _T_279 = s1_tag == cache_tag_s1_entry_r_data; // @[icache.scala 129:23]
  wire  s1_hit = _T_279 & cache_v_s1_entry_r_data; // @[icache.scala 129:40]
  wire  _T_287 = io_in_resp_ready & s1_hit; // @[icache.scala 136:37]
  reg  s1_valid; // @[icache.scala 125:25]
  reg [31:0] _RAND_9;
  wire  _T_288 = ~s1_valid; // @[icache.scala 136:51]
  wire  s0_out_ready = _T_287 | _T_288; // @[icache.scala 136:48]
  wire  s0_out_fire = s0_valid & s0_out_ready; // @[icache.scala 116:30]
  wire  _T_268 = ~s0_valid; // @[icache.scala 117:38]
  wire  _T_271 = ~_T_266; // @[icache.scala 118:19]
  wire  _T_272 = _T_271 & s0_out_fire; // @[icache.scala 118:37]
  wire  _T_273 = flush | _T_272; // @[icache.scala 118:15]
  wire  _T_274 = ~flush; // @[icache.scala 120:15]
  wire  _T_276 = _T_274 & _T_266; // @[icache.scala 120:22]
  wire  _GEN_274 = _T_276 | s0_valid; // @[icache.scala 120:43]
  reg  s1_in_is_cached; // @[Reg.scala 27:20]
  reg [31:0] _RAND_10;
  reg [1:0] s1_in_len; // @[Reg.scala 27:20]
  reg [31:0] _RAND_11;
  reg [3:0] s1_in_strb; // @[Reg.scala 27:20]
  reg [31:0] _RAND_12;
  reg  s1_req; // @[icache.scala 130:23]
  reg [31:0] _RAND_13;
  reg  s1_resp; // @[icache.scala 131:24]
  reg [31:0] _RAND_14;
  wire  _T_280 = s1_req | s1_resp; // @[icache.scala 132:46]
  wire  s1_ex_wait_en = io_ex_flush & _T_280; // @[icache.scala 132:35]
  reg  s1_ex_wait; // @[Reg.scala 27:20]
  reg [31:0] _RAND_15;
  wire  _T_281 = ~s1_req; // @[icache.scala 134:37]
  wire  _T_282 = io_ex_flush & _T_281; // @[icache.scala 134:34]
  wire  _T_283 = ~s1_resp; // @[icache.scala 134:48]
  wire  _T_284 = _T_282 & _T_283; // @[icache.scala 134:45]
  wire  _T_285 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_286 = s1_ex_wait & _T_285; // @[icache.scala 135:17]
  wire  s1_ex_flush = _T_284 | _T_286; // @[icache.scala 134:58]
  wire  _T_290 = s1_valid & s1_hit; // @[icache.scala 137:32]
  wire  _T_291 = ~s1_ex_wait; // @[icache.scala 137:45]
  wire  _T_293 = ~s0_out_fire; // @[icache.scala 139:25]
  wire  _T_294 = io_in_resp_ready & io_in_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_295 = _T_293 & _T_294; // @[icache.scala 139:37]
  wire  _T_296 = s1_ex_flush | _T_295; // @[icache.scala 139:21]
  wire  _T_298 = io_br_flush & _T_294; // @[icache.scala 140:18]
  wire  _T_299 = _T_296 | _T_298; // @[icache.scala 139:59]
  wire  _T_300 = ~s1_ex_flush; // @[icache.scala 142:15]
  wire  _T_301 = _T_300 & s0_out_fire; // @[icache.scala 142:28]
  wire  _GEN_283 = _T_301 | s1_valid; // @[icache.scala 142:43]
  wire  _T_303 = _T & s1_valid; // @[icache.scala 146:22]
  wire  _T_304 = ~s1_hit; // @[icache.scala 146:37]
  wire  _T_305 = _T_303 & _T_304; // @[icache.scala 146:34]
  wire  _T_307 = _T_305 & _T_283; // @[icache.scala 146:45]
  wire  _GEN_285 = _T_307 | s1_req; // @[icache.scala 146:58]
  wire  _T_308 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_309 = s1_req & _T_308; // @[icache.scala 147:16]
  wire  _GEN_287 = _T_309 | s1_resp; // @[icache.scala 147:38]
  wire  _T_311 = s1_resp & _T_285; // @[icache.scala 151:17]
  assign cache_v_s1_entry_r_addr = s1_in_addr[7:0];
  assign cache_v_s1_entry_r_data = cache_v[cache_v_s1_entry_r_addr]; // @[icache.scala 91:18]
  assign cache_v__T_8_data = 1'h0;
  assign cache_v__T_8_addr = _T_6[7:0];
  assign cache_v__T_8_mask = 1'h1;
  assign cache_v__T_8_en = _T_1 & _T_5;
  assign cache_v__T_10_data = 1'h0;
  assign cache_v__T_10_addr = 8'h0;
  assign cache_v__T_10_mask = 1'h1;
  assign cache_v__T_10_en = reset;
  assign cache_v__T_11_data = 1'h0;
  assign cache_v__T_11_addr = 8'h1;
  assign cache_v__T_11_mask = 1'h1;
  assign cache_v__T_11_en = reset;
  assign cache_v__T_12_data = 1'h0;
  assign cache_v__T_12_addr = 8'h2;
  assign cache_v__T_12_mask = 1'h1;
  assign cache_v__T_12_en = reset;
  assign cache_v__T_13_data = 1'h0;
  assign cache_v__T_13_addr = 8'h3;
  assign cache_v__T_13_mask = 1'h1;
  assign cache_v__T_13_en = reset;
  assign cache_v__T_14_data = 1'h0;
  assign cache_v__T_14_addr = 8'h4;
  assign cache_v__T_14_mask = 1'h1;
  assign cache_v__T_14_en = reset;
  assign cache_v__T_15_data = 1'h0;
  assign cache_v__T_15_addr = 8'h5;
  assign cache_v__T_15_mask = 1'h1;
  assign cache_v__T_15_en = reset;
  assign cache_v__T_16_data = 1'h0;
  assign cache_v__T_16_addr = 8'h6;
  assign cache_v__T_16_mask = 1'h1;
  assign cache_v__T_16_en = reset;
  assign cache_v__T_17_data = 1'h0;
  assign cache_v__T_17_addr = 8'h7;
  assign cache_v__T_17_mask = 1'h1;
  assign cache_v__T_17_en = reset;
  assign cache_v__T_18_data = 1'h0;
  assign cache_v__T_18_addr = 8'h8;
  assign cache_v__T_18_mask = 1'h1;
  assign cache_v__T_18_en = reset;
  assign cache_v__T_19_data = 1'h0;
  assign cache_v__T_19_addr = 8'h9;
  assign cache_v__T_19_mask = 1'h1;
  assign cache_v__T_19_en = reset;
  assign cache_v__T_20_data = 1'h0;
  assign cache_v__T_20_addr = 8'ha;
  assign cache_v__T_20_mask = 1'h1;
  assign cache_v__T_20_en = reset;
  assign cache_v__T_21_data = 1'h0;
  assign cache_v__T_21_addr = 8'hb;
  assign cache_v__T_21_mask = 1'h1;
  assign cache_v__T_21_en = reset;
  assign cache_v__T_22_data = 1'h0;
  assign cache_v__T_22_addr = 8'hc;
  assign cache_v__T_22_mask = 1'h1;
  assign cache_v__T_22_en = reset;
  assign cache_v__T_23_data = 1'h0;
  assign cache_v__T_23_addr = 8'hd;
  assign cache_v__T_23_mask = 1'h1;
  assign cache_v__T_23_en = reset;
  assign cache_v__T_24_data = 1'h0;
  assign cache_v__T_24_addr = 8'he;
  assign cache_v__T_24_mask = 1'h1;
  assign cache_v__T_24_en = reset;
  assign cache_v__T_25_data = 1'h0;
  assign cache_v__T_25_addr = 8'hf;
  assign cache_v__T_25_mask = 1'h1;
  assign cache_v__T_25_en = reset;
  assign cache_v__T_26_data = 1'h0;
  assign cache_v__T_26_addr = 8'h10;
  assign cache_v__T_26_mask = 1'h1;
  assign cache_v__T_26_en = reset;
  assign cache_v__T_27_data = 1'h0;
  assign cache_v__T_27_addr = 8'h11;
  assign cache_v__T_27_mask = 1'h1;
  assign cache_v__T_27_en = reset;
  assign cache_v__T_28_data = 1'h0;
  assign cache_v__T_28_addr = 8'h12;
  assign cache_v__T_28_mask = 1'h1;
  assign cache_v__T_28_en = reset;
  assign cache_v__T_29_data = 1'h0;
  assign cache_v__T_29_addr = 8'h13;
  assign cache_v__T_29_mask = 1'h1;
  assign cache_v__T_29_en = reset;
  assign cache_v__T_30_data = 1'h0;
  assign cache_v__T_30_addr = 8'h14;
  assign cache_v__T_30_mask = 1'h1;
  assign cache_v__T_30_en = reset;
  assign cache_v__T_31_data = 1'h0;
  assign cache_v__T_31_addr = 8'h15;
  assign cache_v__T_31_mask = 1'h1;
  assign cache_v__T_31_en = reset;
  assign cache_v__T_32_data = 1'h0;
  assign cache_v__T_32_addr = 8'h16;
  assign cache_v__T_32_mask = 1'h1;
  assign cache_v__T_32_en = reset;
  assign cache_v__T_33_data = 1'h0;
  assign cache_v__T_33_addr = 8'h17;
  assign cache_v__T_33_mask = 1'h1;
  assign cache_v__T_33_en = reset;
  assign cache_v__T_34_data = 1'h0;
  assign cache_v__T_34_addr = 8'h18;
  assign cache_v__T_34_mask = 1'h1;
  assign cache_v__T_34_en = reset;
  assign cache_v__T_35_data = 1'h0;
  assign cache_v__T_35_addr = 8'h19;
  assign cache_v__T_35_mask = 1'h1;
  assign cache_v__T_35_en = reset;
  assign cache_v__T_36_data = 1'h0;
  assign cache_v__T_36_addr = 8'h1a;
  assign cache_v__T_36_mask = 1'h1;
  assign cache_v__T_36_en = reset;
  assign cache_v__T_37_data = 1'h0;
  assign cache_v__T_37_addr = 8'h1b;
  assign cache_v__T_37_mask = 1'h1;
  assign cache_v__T_37_en = reset;
  assign cache_v__T_38_data = 1'h0;
  assign cache_v__T_38_addr = 8'h1c;
  assign cache_v__T_38_mask = 1'h1;
  assign cache_v__T_38_en = reset;
  assign cache_v__T_39_data = 1'h0;
  assign cache_v__T_39_addr = 8'h1d;
  assign cache_v__T_39_mask = 1'h1;
  assign cache_v__T_39_en = reset;
  assign cache_v__T_40_data = 1'h0;
  assign cache_v__T_40_addr = 8'h1e;
  assign cache_v__T_40_mask = 1'h1;
  assign cache_v__T_40_en = reset;
  assign cache_v__T_41_data = 1'h0;
  assign cache_v__T_41_addr = 8'h1f;
  assign cache_v__T_41_mask = 1'h1;
  assign cache_v__T_41_en = reset;
  assign cache_v__T_42_data = 1'h0;
  assign cache_v__T_42_addr = 8'h20;
  assign cache_v__T_42_mask = 1'h1;
  assign cache_v__T_42_en = reset;
  assign cache_v__T_43_data = 1'h0;
  assign cache_v__T_43_addr = 8'h21;
  assign cache_v__T_43_mask = 1'h1;
  assign cache_v__T_43_en = reset;
  assign cache_v__T_44_data = 1'h0;
  assign cache_v__T_44_addr = 8'h22;
  assign cache_v__T_44_mask = 1'h1;
  assign cache_v__T_44_en = reset;
  assign cache_v__T_45_data = 1'h0;
  assign cache_v__T_45_addr = 8'h23;
  assign cache_v__T_45_mask = 1'h1;
  assign cache_v__T_45_en = reset;
  assign cache_v__T_46_data = 1'h0;
  assign cache_v__T_46_addr = 8'h24;
  assign cache_v__T_46_mask = 1'h1;
  assign cache_v__T_46_en = reset;
  assign cache_v__T_47_data = 1'h0;
  assign cache_v__T_47_addr = 8'h25;
  assign cache_v__T_47_mask = 1'h1;
  assign cache_v__T_47_en = reset;
  assign cache_v__T_48_data = 1'h0;
  assign cache_v__T_48_addr = 8'h26;
  assign cache_v__T_48_mask = 1'h1;
  assign cache_v__T_48_en = reset;
  assign cache_v__T_49_data = 1'h0;
  assign cache_v__T_49_addr = 8'h27;
  assign cache_v__T_49_mask = 1'h1;
  assign cache_v__T_49_en = reset;
  assign cache_v__T_50_data = 1'h0;
  assign cache_v__T_50_addr = 8'h28;
  assign cache_v__T_50_mask = 1'h1;
  assign cache_v__T_50_en = reset;
  assign cache_v__T_51_data = 1'h0;
  assign cache_v__T_51_addr = 8'h29;
  assign cache_v__T_51_mask = 1'h1;
  assign cache_v__T_51_en = reset;
  assign cache_v__T_52_data = 1'h0;
  assign cache_v__T_52_addr = 8'h2a;
  assign cache_v__T_52_mask = 1'h1;
  assign cache_v__T_52_en = reset;
  assign cache_v__T_53_data = 1'h0;
  assign cache_v__T_53_addr = 8'h2b;
  assign cache_v__T_53_mask = 1'h1;
  assign cache_v__T_53_en = reset;
  assign cache_v__T_54_data = 1'h0;
  assign cache_v__T_54_addr = 8'h2c;
  assign cache_v__T_54_mask = 1'h1;
  assign cache_v__T_54_en = reset;
  assign cache_v__T_55_data = 1'h0;
  assign cache_v__T_55_addr = 8'h2d;
  assign cache_v__T_55_mask = 1'h1;
  assign cache_v__T_55_en = reset;
  assign cache_v__T_56_data = 1'h0;
  assign cache_v__T_56_addr = 8'h2e;
  assign cache_v__T_56_mask = 1'h1;
  assign cache_v__T_56_en = reset;
  assign cache_v__T_57_data = 1'h0;
  assign cache_v__T_57_addr = 8'h2f;
  assign cache_v__T_57_mask = 1'h1;
  assign cache_v__T_57_en = reset;
  assign cache_v__T_58_data = 1'h0;
  assign cache_v__T_58_addr = 8'h30;
  assign cache_v__T_58_mask = 1'h1;
  assign cache_v__T_58_en = reset;
  assign cache_v__T_59_data = 1'h0;
  assign cache_v__T_59_addr = 8'h31;
  assign cache_v__T_59_mask = 1'h1;
  assign cache_v__T_59_en = reset;
  assign cache_v__T_60_data = 1'h0;
  assign cache_v__T_60_addr = 8'h32;
  assign cache_v__T_60_mask = 1'h1;
  assign cache_v__T_60_en = reset;
  assign cache_v__T_61_data = 1'h0;
  assign cache_v__T_61_addr = 8'h33;
  assign cache_v__T_61_mask = 1'h1;
  assign cache_v__T_61_en = reset;
  assign cache_v__T_62_data = 1'h0;
  assign cache_v__T_62_addr = 8'h34;
  assign cache_v__T_62_mask = 1'h1;
  assign cache_v__T_62_en = reset;
  assign cache_v__T_63_data = 1'h0;
  assign cache_v__T_63_addr = 8'h35;
  assign cache_v__T_63_mask = 1'h1;
  assign cache_v__T_63_en = reset;
  assign cache_v__T_64_data = 1'h0;
  assign cache_v__T_64_addr = 8'h36;
  assign cache_v__T_64_mask = 1'h1;
  assign cache_v__T_64_en = reset;
  assign cache_v__T_65_data = 1'h0;
  assign cache_v__T_65_addr = 8'h37;
  assign cache_v__T_65_mask = 1'h1;
  assign cache_v__T_65_en = reset;
  assign cache_v__T_66_data = 1'h0;
  assign cache_v__T_66_addr = 8'h38;
  assign cache_v__T_66_mask = 1'h1;
  assign cache_v__T_66_en = reset;
  assign cache_v__T_67_data = 1'h0;
  assign cache_v__T_67_addr = 8'h39;
  assign cache_v__T_67_mask = 1'h1;
  assign cache_v__T_67_en = reset;
  assign cache_v__T_68_data = 1'h0;
  assign cache_v__T_68_addr = 8'h3a;
  assign cache_v__T_68_mask = 1'h1;
  assign cache_v__T_68_en = reset;
  assign cache_v__T_69_data = 1'h0;
  assign cache_v__T_69_addr = 8'h3b;
  assign cache_v__T_69_mask = 1'h1;
  assign cache_v__T_69_en = reset;
  assign cache_v__T_70_data = 1'h0;
  assign cache_v__T_70_addr = 8'h3c;
  assign cache_v__T_70_mask = 1'h1;
  assign cache_v__T_70_en = reset;
  assign cache_v__T_71_data = 1'h0;
  assign cache_v__T_71_addr = 8'h3d;
  assign cache_v__T_71_mask = 1'h1;
  assign cache_v__T_71_en = reset;
  assign cache_v__T_72_data = 1'h0;
  assign cache_v__T_72_addr = 8'h3e;
  assign cache_v__T_72_mask = 1'h1;
  assign cache_v__T_72_en = reset;
  assign cache_v__T_73_data = 1'h0;
  assign cache_v__T_73_addr = 8'h3f;
  assign cache_v__T_73_mask = 1'h1;
  assign cache_v__T_73_en = reset;
  assign cache_v__T_74_data = 1'h0;
  assign cache_v__T_74_addr = 8'h40;
  assign cache_v__T_74_mask = 1'h1;
  assign cache_v__T_74_en = reset;
  assign cache_v__T_75_data = 1'h0;
  assign cache_v__T_75_addr = 8'h41;
  assign cache_v__T_75_mask = 1'h1;
  assign cache_v__T_75_en = reset;
  assign cache_v__T_76_data = 1'h0;
  assign cache_v__T_76_addr = 8'h42;
  assign cache_v__T_76_mask = 1'h1;
  assign cache_v__T_76_en = reset;
  assign cache_v__T_77_data = 1'h0;
  assign cache_v__T_77_addr = 8'h43;
  assign cache_v__T_77_mask = 1'h1;
  assign cache_v__T_77_en = reset;
  assign cache_v__T_78_data = 1'h0;
  assign cache_v__T_78_addr = 8'h44;
  assign cache_v__T_78_mask = 1'h1;
  assign cache_v__T_78_en = reset;
  assign cache_v__T_79_data = 1'h0;
  assign cache_v__T_79_addr = 8'h45;
  assign cache_v__T_79_mask = 1'h1;
  assign cache_v__T_79_en = reset;
  assign cache_v__T_80_data = 1'h0;
  assign cache_v__T_80_addr = 8'h46;
  assign cache_v__T_80_mask = 1'h1;
  assign cache_v__T_80_en = reset;
  assign cache_v__T_81_data = 1'h0;
  assign cache_v__T_81_addr = 8'h47;
  assign cache_v__T_81_mask = 1'h1;
  assign cache_v__T_81_en = reset;
  assign cache_v__T_82_data = 1'h0;
  assign cache_v__T_82_addr = 8'h48;
  assign cache_v__T_82_mask = 1'h1;
  assign cache_v__T_82_en = reset;
  assign cache_v__T_83_data = 1'h0;
  assign cache_v__T_83_addr = 8'h49;
  assign cache_v__T_83_mask = 1'h1;
  assign cache_v__T_83_en = reset;
  assign cache_v__T_84_data = 1'h0;
  assign cache_v__T_84_addr = 8'h4a;
  assign cache_v__T_84_mask = 1'h1;
  assign cache_v__T_84_en = reset;
  assign cache_v__T_85_data = 1'h0;
  assign cache_v__T_85_addr = 8'h4b;
  assign cache_v__T_85_mask = 1'h1;
  assign cache_v__T_85_en = reset;
  assign cache_v__T_86_data = 1'h0;
  assign cache_v__T_86_addr = 8'h4c;
  assign cache_v__T_86_mask = 1'h1;
  assign cache_v__T_86_en = reset;
  assign cache_v__T_87_data = 1'h0;
  assign cache_v__T_87_addr = 8'h4d;
  assign cache_v__T_87_mask = 1'h1;
  assign cache_v__T_87_en = reset;
  assign cache_v__T_88_data = 1'h0;
  assign cache_v__T_88_addr = 8'h4e;
  assign cache_v__T_88_mask = 1'h1;
  assign cache_v__T_88_en = reset;
  assign cache_v__T_89_data = 1'h0;
  assign cache_v__T_89_addr = 8'h4f;
  assign cache_v__T_89_mask = 1'h1;
  assign cache_v__T_89_en = reset;
  assign cache_v__T_90_data = 1'h0;
  assign cache_v__T_90_addr = 8'h50;
  assign cache_v__T_90_mask = 1'h1;
  assign cache_v__T_90_en = reset;
  assign cache_v__T_91_data = 1'h0;
  assign cache_v__T_91_addr = 8'h51;
  assign cache_v__T_91_mask = 1'h1;
  assign cache_v__T_91_en = reset;
  assign cache_v__T_92_data = 1'h0;
  assign cache_v__T_92_addr = 8'h52;
  assign cache_v__T_92_mask = 1'h1;
  assign cache_v__T_92_en = reset;
  assign cache_v__T_93_data = 1'h0;
  assign cache_v__T_93_addr = 8'h53;
  assign cache_v__T_93_mask = 1'h1;
  assign cache_v__T_93_en = reset;
  assign cache_v__T_94_data = 1'h0;
  assign cache_v__T_94_addr = 8'h54;
  assign cache_v__T_94_mask = 1'h1;
  assign cache_v__T_94_en = reset;
  assign cache_v__T_95_data = 1'h0;
  assign cache_v__T_95_addr = 8'h55;
  assign cache_v__T_95_mask = 1'h1;
  assign cache_v__T_95_en = reset;
  assign cache_v__T_96_data = 1'h0;
  assign cache_v__T_96_addr = 8'h56;
  assign cache_v__T_96_mask = 1'h1;
  assign cache_v__T_96_en = reset;
  assign cache_v__T_97_data = 1'h0;
  assign cache_v__T_97_addr = 8'h57;
  assign cache_v__T_97_mask = 1'h1;
  assign cache_v__T_97_en = reset;
  assign cache_v__T_98_data = 1'h0;
  assign cache_v__T_98_addr = 8'h58;
  assign cache_v__T_98_mask = 1'h1;
  assign cache_v__T_98_en = reset;
  assign cache_v__T_99_data = 1'h0;
  assign cache_v__T_99_addr = 8'h59;
  assign cache_v__T_99_mask = 1'h1;
  assign cache_v__T_99_en = reset;
  assign cache_v__T_100_data = 1'h0;
  assign cache_v__T_100_addr = 8'h5a;
  assign cache_v__T_100_mask = 1'h1;
  assign cache_v__T_100_en = reset;
  assign cache_v__T_101_data = 1'h0;
  assign cache_v__T_101_addr = 8'h5b;
  assign cache_v__T_101_mask = 1'h1;
  assign cache_v__T_101_en = reset;
  assign cache_v__T_102_data = 1'h0;
  assign cache_v__T_102_addr = 8'h5c;
  assign cache_v__T_102_mask = 1'h1;
  assign cache_v__T_102_en = reset;
  assign cache_v__T_103_data = 1'h0;
  assign cache_v__T_103_addr = 8'h5d;
  assign cache_v__T_103_mask = 1'h1;
  assign cache_v__T_103_en = reset;
  assign cache_v__T_104_data = 1'h0;
  assign cache_v__T_104_addr = 8'h5e;
  assign cache_v__T_104_mask = 1'h1;
  assign cache_v__T_104_en = reset;
  assign cache_v__T_105_data = 1'h0;
  assign cache_v__T_105_addr = 8'h5f;
  assign cache_v__T_105_mask = 1'h1;
  assign cache_v__T_105_en = reset;
  assign cache_v__T_106_data = 1'h0;
  assign cache_v__T_106_addr = 8'h60;
  assign cache_v__T_106_mask = 1'h1;
  assign cache_v__T_106_en = reset;
  assign cache_v__T_107_data = 1'h0;
  assign cache_v__T_107_addr = 8'h61;
  assign cache_v__T_107_mask = 1'h1;
  assign cache_v__T_107_en = reset;
  assign cache_v__T_108_data = 1'h0;
  assign cache_v__T_108_addr = 8'h62;
  assign cache_v__T_108_mask = 1'h1;
  assign cache_v__T_108_en = reset;
  assign cache_v__T_109_data = 1'h0;
  assign cache_v__T_109_addr = 8'h63;
  assign cache_v__T_109_mask = 1'h1;
  assign cache_v__T_109_en = reset;
  assign cache_v__T_110_data = 1'h0;
  assign cache_v__T_110_addr = 8'h64;
  assign cache_v__T_110_mask = 1'h1;
  assign cache_v__T_110_en = reset;
  assign cache_v__T_111_data = 1'h0;
  assign cache_v__T_111_addr = 8'h65;
  assign cache_v__T_111_mask = 1'h1;
  assign cache_v__T_111_en = reset;
  assign cache_v__T_112_data = 1'h0;
  assign cache_v__T_112_addr = 8'h66;
  assign cache_v__T_112_mask = 1'h1;
  assign cache_v__T_112_en = reset;
  assign cache_v__T_113_data = 1'h0;
  assign cache_v__T_113_addr = 8'h67;
  assign cache_v__T_113_mask = 1'h1;
  assign cache_v__T_113_en = reset;
  assign cache_v__T_114_data = 1'h0;
  assign cache_v__T_114_addr = 8'h68;
  assign cache_v__T_114_mask = 1'h1;
  assign cache_v__T_114_en = reset;
  assign cache_v__T_115_data = 1'h0;
  assign cache_v__T_115_addr = 8'h69;
  assign cache_v__T_115_mask = 1'h1;
  assign cache_v__T_115_en = reset;
  assign cache_v__T_116_data = 1'h0;
  assign cache_v__T_116_addr = 8'h6a;
  assign cache_v__T_116_mask = 1'h1;
  assign cache_v__T_116_en = reset;
  assign cache_v__T_117_data = 1'h0;
  assign cache_v__T_117_addr = 8'h6b;
  assign cache_v__T_117_mask = 1'h1;
  assign cache_v__T_117_en = reset;
  assign cache_v__T_118_data = 1'h0;
  assign cache_v__T_118_addr = 8'h6c;
  assign cache_v__T_118_mask = 1'h1;
  assign cache_v__T_118_en = reset;
  assign cache_v__T_119_data = 1'h0;
  assign cache_v__T_119_addr = 8'h6d;
  assign cache_v__T_119_mask = 1'h1;
  assign cache_v__T_119_en = reset;
  assign cache_v__T_120_data = 1'h0;
  assign cache_v__T_120_addr = 8'h6e;
  assign cache_v__T_120_mask = 1'h1;
  assign cache_v__T_120_en = reset;
  assign cache_v__T_121_data = 1'h0;
  assign cache_v__T_121_addr = 8'h6f;
  assign cache_v__T_121_mask = 1'h1;
  assign cache_v__T_121_en = reset;
  assign cache_v__T_122_data = 1'h0;
  assign cache_v__T_122_addr = 8'h70;
  assign cache_v__T_122_mask = 1'h1;
  assign cache_v__T_122_en = reset;
  assign cache_v__T_123_data = 1'h0;
  assign cache_v__T_123_addr = 8'h71;
  assign cache_v__T_123_mask = 1'h1;
  assign cache_v__T_123_en = reset;
  assign cache_v__T_124_data = 1'h0;
  assign cache_v__T_124_addr = 8'h72;
  assign cache_v__T_124_mask = 1'h1;
  assign cache_v__T_124_en = reset;
  assign cache_v__T_125_data = 1'h0;
  assign cache_v__T_125_addr = 8'h73;
  assign cache_v__T_125_mask = 1'h1;
  assign cache_v__T_125_en = reset;
  assign cache_v__T_126_data = 1'h0;
  assign cache_v__T_126_addr = 8'h74;
  assign cache_v__T_126_mask = 1'h1;
  assign cache_v__T_126_en = reset;
  assign cache_v__T_127_data = 1'h0;
  assign cache_v__T_127_addr = 8'h75;
  assign cache_v__T_127_mask = 1'h1;
  assign cache_v__T_127_en = reset;
  assign cache_v__T_128_data = 1'h0;
  assign cache_v__T_128_addr = 8'h76;
  assign cache_v__T_128_mask = 1'h1;
  assign cache_v__T_128_en = reset;
  assign cache_v__T_129_data = 1'h0;
  assign cache_v__T_129_addr = 8'h77;
  assign cache_v__T_129_mask = 1'h1;
  assign cache_v__T_129_en = reset;
  assign cache_v__T_130_data = 1'h0;
  assign cache_v__T_130_addr = 8'h78;
  assign cache_v__T_130_mask = 1'h1;
  assign cache_v__T_130_en = reset;
  assign cache_v__T_131_data = 1'h0;
  assign cache_v__T_131_addr = 8'h79;
  assign cache_v__T_131_mask = 1'h1;
  assign cache_v__T_131_en = reset;
  assign cache_v__T_132_data = 1'h0;
  assign cache_v__T_132_addr = 8'h7a;
  assign cache_v__T_132_mask = 1'h1;
  assign cache_v__T_132_en = reset;
  assign cache_v__T_133_data = 1'h0;
  assign cache_v__T_133_addr = 8'h7b;
  assign cache_v__T_133_mask = 1'h1;
  assign cache_v__T_133_en = reset;
  assign cache_v__T_134_data = 1'h0;
  assign cache_v__T_134_addr = 8'h7c;
  assign cache_v__T_134_mask = 1'h1;
  assign cache_v__T_134_en = reset;
  assign cache_v__T_135_data = 1'h0;
  assign cache_v__T_135_addr = 8'h7d;
  assign cache_v__T_135_mask = 1'h1;
  assign cache_v__T_135_en = reset;
  assign cache_v__T_136_data = 1'h0;
  assign cache_v__T_136_addr = 8'h7e;
  assign cache_v__T_136_mask = 1'h1;
  assign cache_v__T_136_en = reset;
  assign cache_v__T_137_data = 1'h0;
  assign cache_v__T_137_addr = 8'h7f;
  assign cache_v__T_137_mask = 1'h1;
  assign cache_v__T_137_en = reset;
  assign cache_v__T_138_data = 1'h0;
  assign cache_v__T_138_addr = 8'h80;
  assign cache_v__T_138_mask = 1'h1;
  assign cache_v__T_138_en = reset;
  assign cache_v__T_139_data = 1'h0;
  assign cache_v__T_139_addr = 8'h81;
  assign cache_v__T_139_mask = 1'h1;
  assign cache_v__T_139_en = reset;
  assign cache_v__T_140_data = 1'h0;
  assign cache_v__T_140_addr = 8'h82;
  assign cache_v__T_140_mask = 1'h1;
  assign cache_v__T_140_en = reset;
  assign cache_v__T_141_data = 1'h0;
  assign cache_v__T_141_addr = 8'h83;
  assign cache_v__T_141_mask = 1'h1;
  assign cache_v__T_141_en = reset;
  assign cache_v__T_142_data = 1'h0;
  assign cache_v__T_142_addr = 8'h84;
  assign cache_v__T_142_mask = 1'h1;
  assign cache_v__T_142_en = reset;
  assign cache_v__T_143_data = 1'h0;
  assign cache_v__T_143_addr = 8'h85;
  assign cache_v__T_143_mask = 1'h1;
  assign cache_v__T_143_en = reset;
  assign cache_v__T_144_data = 1'h0;
  assign cache_v__T_144_addr = 8'h86;
  assign cache_v__T_144_mask = 1'h1;
  assign cache_v__T_144_en = reset;
  assign cache_v__T_145_data = 1'h0;
  assign cache_v__T_145_addr = 8'h87;
  assign cache_v__T_145_mask = 1'h1;
  assign cache_v__T_145_en = reset;
  assign cache_v__T_146_data = 1'h0;
  assign cache_v__T_146_addr = 8'h88;
  assign cache_v__T_146_mask = 1'h1;
  assign cache_v__T_146_en = reset;
  assign cache_v__T_147_data = 1'h0;
  assign cache_v__T_147_addr = 8'h89;
  assign cache_v__T_147_mask = 1'h1;
  assign cache_v__T_147_en = reset;
  assign cache_v__T_148_data = 1'h0;
  assign cache_v__T_148_addr = 8'h8a;
  assign cache_v__T_148_mask = 1'h1;
  assign cache_v__T_148_en = reset;
  assign cache_v__T_149_data = 1'h0;
  assign cache_v__T_149_addr = 8'h8b;
  assign cache_v__T_149_mask = 1'h1;
  assign cache_v__T_149_en = reset;
  assign cache_v__T_150_data = 1'h0;
  assign cache_v__T_150_addr = 8'h8c;
  assign cache_v__T_150_mask = 1'h1;
  assign cache_v__T_150_en = reset;
  assign cache_v__T_151_data = 1'h0;
  assign cache_v__T_151_addr = 8'h8d;
  assign cache_v__T_151_mask = 1'h1;
  assign cache_v__T_151_en = reset;
  assign cache_v__T_152_data = 1'h0;
  assign cache_v__T_152_addr = 8'h8e;
  assign cache_v__T_152_mask = 1'h1;
  assign cache_v__T_152_en = reset;
  assign cache_v__T_153_data = 1'h0;
  assign cache_v__T_153_addr = 8'h8f;
  assign cache_v__T_153_mask = 1'h1;
  assign cache_v__T_153_en = reset;
  assign cache_v__T_154_data = 1'h0;
  assign cache_v__T_154_addr = 8'h90;
  assign cache_v__T_154_mask = 1'h1;
  assign cache_v__T_154_en = reset;
  assign cache_v__T_155_data = 1'h0;
  assign cache_v__T_155_addr = 8'h91;
  assign cache_v__T_155_mask = 1'h1;
  assign cache_v__T_155_en = reset;
  assign cache_v__T_156_data = 1'h0;
  assign cache_v__T_156_addr = 8'h92;
  assign cache_v__T_156_mask = 1'h1;
  assign cache_v__T_156_en = reset;
  assign cache_v__T_157_data = 1'h0;
  assign cache_v__T_157_addr = 8'h93;
  assign cache_v__T_157_mask = 1'h1;
  assign cache_v__T_157_en = reset;
  assign cache_v__T_158_data = 1'h0;
  assign cache_v__T_158_addr = 8'h94;
  assign cache_v__T_158_mask = 1'h1;
  assign cache_v__T_158_en = reset;
  assign cache_v__T_159_data = 1'h0;
  assign cache_v__T_159_addr = 8'h95;
  assign cache_v__T_159_mask = 1'h1;
  assign cache_v__T_159_en = reset;
  assign cache_v__T_160_data = 1'h0;
  assign cache_v__T_160_addr = 8'h96;
  assign cache_v__T_160_mask = 1'h1;
  assign cache_v__T_160_en = reset;
  assign cache_v__T_161_data = 1'h0;
  assign cache_v__T_161_addr = 8'h97;
  assign cache_v__T_161_mask = 1'h1;
  assign cache_v__T_161_en = reset;
  assign cache_v__T_162_data = 1'h0;
  assign cache_v__T_162_addr = 8'h98;
  assign cache_v__T_162_mask = 1'h1;
  assign cache_v__T_162_en = reset;
  assign cache_v__T_163_data = 1'h0;
  assign cache_v__T_163_addr = 8'h99;
  assign cache_v__T_163_mask = 1'h1;
  assign cache_v__T_163_en = reset;
  assign cache_v__T_164_data = 1'h0;
  assign cache_v__T_164_addr = 8'h9a;
  assign cache_v__T_164_mask = 1'h1;
  assign cache_v__T_164_en = reset;
  assign cache_v__T_165_data = 1'h0;
  assign cache_v__T_165_addr = 8'h9b;
  assign cache_v__T_165_mask = 1'h1;
  assign cache_v__T_165_en = reset;
  assign cache_v__T_166_data = 1'h0;
  assign cache_v__T_166_addr = 8'h9c;
  assign cache_v__T_166_mask = 1'h1;
  assign cache_v__T_166_en = reset;
  assign cache_v__T_167_data = 1'h0;
  assign cache_v__T_167_addr = 8'h9d;
  assign cache_v__T_167_mask = 1'h1;
  assign cache_v__T_167_en = reset;
  assign cache_v__T_168_data = 1'h0;
  assign cache_v__T_168_addr = 8'h9e;
  assign cache_v__T_168_mask = 1'h1;
  assign cache_v__T_168_en = reset;
  assign cache_v__T_169_data = 1'h0;
  assign cache_v__T_169_addr = 8'h9f;
  assign cache_v__T_169_mask = 1'h1;
  assign cache_v__T_169_en = reset;
  assign cache_v__T_170_data = 1'h0;
  assign cache_v__T_170_addr = 8'ha0;
  assign cache_v__T_170_mask = 1'h1;
  assign cache_v__T_170_en = reset;
  assign cache_v__T_171_data = 1'h0;
  assign cache_v__T_171_addr = 8'ha1;
  assign cache_v__T_171_mask = 1'h1;
  assign cache_v__T_171_en = reset;
  assign cache_v__T_172_data = 1'h0;
  assign cache_v__T_172_addr = 8'ha2;
  assign cache_v__T_172_mask = 1'h1;
  assign cache_v__T_172_en = reset;
  assign cache_v__T_173_data = 1'h0;
  assign cache_v__T_173_addr = 8'ha3;
  assign cache_v__T_173_mask = 1'h1;
  assign cache_v__T_173_en = reset;
  assign cache_v__T_174_data = 1'h0;
  assign cache_v__T_174_addr = 8'ha4;
  assign cache_v__T_174_mask = 1'h1;
  assign cache_v__T_174_en = reset;
  assign cache_v__T_175_data = 1'h0;
  assign cache_v__T_175_addr = 8'ha5;
  assign cache_v__T_175_mask = 1'h1;
  assign cache_v__T_175_en = reset;
  assign cache_v__T_176_data = 1'h0;
  assign cache_v__T_176_addr = 8'ha6;
  assign cache_v__T_176_mask = 1'h1;
  assign cache_v__T_176_en = reset;
  assign cache_v__T_177_data = 1'h0;
  assign cache_v__T_177_addr = 8'ha7;
  assign cache_v__T_177_mask = 1'h1;
  assign cache_v__T_177_en = reset;
  assign cache_v__T_178_data = 1'h0;
  assign cache_v__T_178_addr = 8'ha8;
  assign cache_v__T_178_mask = 1'h1;
  assign cache_v__T_178_en = reset;
  assign cache_v__T_179_data = 1'h0;
  assign cache_v__T_179_addr = 8'ha9;
  assign cache_v__T_179_mask = 1'h1;
  assign cache_v__T_179_en = reset;
  assign cache_v__T_180_data = 1'h0;
  assign cache_v__T_180_addr = 8'haa;
  assign cache_v__T_180_mask = 1'h1;
  assign cache_v__T_180_en = reset;
  assign cache_v__T_181_data = 1'h0;
  assign cache_v__T_181_addr = 8'hab;
  assign cache_v__T_181_mask = 1'h1;
  assign cache_v__T_181_en = reset;
  assign cache_v__T_182_data = 1'h0;
  assign cache_v__T_182_addr = 8'hac;
  assign cache_v__T_182_mask = 1'h1;
  assign cache_v__T_182_en = reset;
  assign cache_v__T_183_data = 1'h0;
  assign cache_v__T_183_addr = 8'had;
  assign cache_v__T_183_mask = 1'h1;
  assign cache_v__T_183_en = reset;
  assign cache_v__T_184_data = 1'h0;
  assign cache_v__T_184_addr = 8'hae;
  assign cache_v__T_184_mask = 1'h1;
  assign cache_v__T_184_en = reset;
  assign cache_v__T_185_data = 1'h0;
  assign cache_v__T_185_addr = 8'haf;
  assign cache_v__T_185_mask = 1'h1;
  assign cache_v__T_185_en = reset;
  assign cache_v__T_186_data = 1'h0;
  assign cache_v__T_186_addr = 8'hb0;
  assign cache_v__T_186_mask = 1'h1;
  assign cache_v__T_186_en = reset;
  assign cache_v__T_187_data = 1'h0;
  assign cache_v__T_187_addr = 8'hb1;
  assign cache_v__T_187_mask = 1'h1;
  assign cache_v__T_187_en = reset;
  assign cache_v__T_188_data = 1'h0;
  assign cache_v__T_188_addr = 8'hb2;
  assign cache_v__T_188_mask = 1'h1;
  assign cache_v__T_188_en = reset;
  assign cache_v__T_189_data = 1'h0;
  assign cache_v__T_189_addr = 8'hb3;
  assign cache_v__T_189_mask = 1'h1;
  assign cache_v__T_189_en = reset;
  assign cache_v__T_190_data = 1'h0;
  assign cache_v__T_190_addr = 8'hb4;
  assign cache_v__T_190_mask = 1'h1;
  assign cache_v__T_190_en = reset;
  assign cache_v__T_191_data = 1'h0;
  assign cache_v__T_191_addr = 8'hb5;
  assign cache_v__T_191_mask = 1'h1;
  assign cache_v__T_191_en = reset;
  assign cache_v__T_192_data = 1'h0;
  assign cache_v__T_192_addr = 8'hb6;
  assign cache_v__T_192_mask = 1'h1;
  assign cache_v__T_192_en = reset;
  assign cache_v__T_193_data = 1'h0;
  assign cache_v__T_193_addr = 8'hb7;
  assign cache_v__T_193_mask = 1'h1;
  assign cache_v__T_193_en = reset;
  assign cache_v__T_194_data = 1'h0;
  assign cache_v__T_194_addr = 8'hb8;
  assign cache_v__T_194_mask = 1'h1;
  assign cache_v__T_194_en = reset;
  assign cache_v__T_195_data = 1'h0;
  assign cache_v__T_195_addr = 8'hb9;
  assign cache_v__T_195_mask = 1'h1;
  assign cache_v__T_195_en = reset;
  assign cache_v__T_196_data = 1'h0;
  assign cache_v__T_196_addr = 8'hba;
  assign cache_v__T_196_mask = 1'h1;
  assign cache_v__T_196_en = reset;
  assign cache_v__T_197_data = 1'h0;
  assign cache_v__T_197_addr = 8'hbb;
  assign cache_v__T_197_mask = 1'h1;
  assign cache_v__T_197_en = reset;
  assign cache_v__T_198_data = 1'h0;
  assign cache_v__T_198_addr = 8'hbc;
  assign cache_v__T_198_mask = 1'h1;
  assign cache_v__T_198_en = reset;
  assign cache_v__T_199_data = 1'h0;
  assign cache_v__T_199_addr = 8'hbd;
  assign cache_v__T_199_mask = 1'h1;
  assign cache_v__T_199_en = reset;
  assign cache_v__T_200_data = 1'h0;
  assign cache_v__T_200_addr = 8'hbe;
  assign cache_v__T_200_mask = 1'h1;
  assign cache_v__T_200_en = reset;
  assign cache_v__T_201_data = 1'h0;
  assign cache_v__T_201_addr = 8'hbf;
  assign cache_v__T_201_mask = 1'h1;
  assign cache_v__T_201_en = reset;
  assign cache_v__T_202_data = 1'h0;
  assign cache_v__T_202_addr = 8'hc0;
  assign cache_v__T_202_mask = 1'h1;
  assign cache_v__T_202_en = reset;
  assign cache_v__T_203_data = 1'h0;
  assign cache_v__T_203_addr = 8'hc1;
  assign cache_v__T_203_mask = 1'h1;
  assign cache_v__T_203_en = reset;
  assign cache_v__T_204_data = 1'h0;
  assign cache_v__T_204_addr = 8'hc2;
  assign cache_v__T_204_mask = 1'h1;
  assign cache_v__T_204_en = reset;
  assign cache_v__T_205_data = 1'h0;
  assign cache_v__T_205_addr = 8'hc3;
  assign cache_v__T_205_mask = 1'h1;
  assign cache_v__T_205_en = reset;
  assign cache_v__T_206_data = 1'h0;
  assign cache_v__T_206_addr = 8'hc4;
  assign cache_v__T_206_mask = 1'h1;
  assign cache_v__T_206_en = reset;
  assign cache_v__T_207_data = 1'h0;
  assign cache_v__T_207_addr = 8'hc5;
  assign cache_v__T_207_mask = 1'h1;
  assign cache_v__T_207_en = reset;
  assign cache_v__T_208_data = 1'h0;
  assign cache_v__T_208_addr = 8'hc6;
  assign cache_v__T_208_mask = 1'h1;
  assign cache_v__T_208_en = reset;
  assign cache_v__T_209_data = 1'h0;
  assign cache_v__T_209_addr = 8'hc7;
  assign cache_v__T_209_mask = 1'h1;
  assign cache_v__T_209_en = reset;
  assign cache_v__T_210_data = 1'h0;
  assign cache_v__T_210_addr = 8'hc8;
  assign cache_v__T_210_mask = 1'h1;
  assign cache_v__T_210_en = reset;
  assign cache_v__T_211_data = 1'h0;
  assign cache_v__T_211_addr = 8'hc9;
  assign cache_v__T_211_mask = 1'h1;
  assign cache_v__T_211_en = reset;
  assign cache_v__T_212_data = 1'h0;
  assign cache_v__T_212_addr = 8'hca;
  assign cache_v__T_212_mask = 1'h1;
  assign cache_v__T_212_en = reset;
  assign cache_v__T_213_data = 1'h0;
  assign cache_v__T_213_addr = 8'hcb;
  assign cache_v__T_213_mask = 1'h1;
  assign cache_v__T_213_en = reset;
  assign cache_v__T_214_data = 1'h0;
  assign cache_v__T_214_addr = 8'hcc;
  assign cache_v__T_214_mask = 1'h1;
  assign cache_v__T_214_en = reset;
  assign cache_v__T_215_data = 1'h0;
  assign cache_v__T_215_addr = 8'hcd;
  assign cache_v__T_215_mask = 1'h1;
  assign cache_v__T_215_en = reset;
  assign cache_v__T_216_data = 1'h0;
  assign cache_v__T_216_addr = 8'hce;
  assign cache_v__T_216_mask = 1'h1;
  assign cache_v__T_216_en = reset;
  assign cache_v__T_217_data = 1'h0;
  assign cache_v__T_217_addr = 8'hcf;
  assign cache_v__T_217_mask = 1'h1;
  assign cache_v__T_217_en = reset;
  assign cache_v__T_218_data = 1'h0;
  assign cache_v__T_218_addr = 8'hd0;
  assign cache_v__T_218_mask = 1'h1;
  assign cache_v__T_218_en = reset;
  assign cache_v__T_219_data = 1'h0;
  assign cache_v__T_219_addr = 8'hd1;
  assign cache_v__T_219_mask = 1'h1;
  assign cache_v__T_219_en = reset;
  assign cache_v__T_220_data = 1'h0;
  assign cache_v__T_220_addr = 8'hd2;
  assign cache_v__T_220_mask = 1'h1;
  assign cache_v__T_220_en = reset;
  assign cache_v__T_221_data = 1'h0;
  assign cache_v__T_221_addr = 8'hd3;
  assign cache_v__T_221_mask = 1'h1;
  assign cache_v__T_221_en = reset;
  assign cache_v__T_222_data = 1'h0;
  assign cache_v__T_222_addr = 8'hd4;
  assign cache_v__T_222_mask = 1'h1;
  assign cache_v__T_222_en = reset;
  assign cache_v__T_223_data = 1'h0;
  assign cache_v__T_223_addr = 8'hd5;
  assign cache_v__T_223_mask = 1'h1;
  assign cache_v__T_223_en = reset;
  assign cache_v__T_224_data = 1'h0;
  assign cache_v__T_224_addr = 8'hd6;
  assign cache_v__T_224_mask = 1'h1;
  assign cache_v__T_224_en = reset;
  assign cache_v__T_225_data = 1'h0;
  assign cache_v__T_225_addr = 8'hd7;
  assign cache_v__T_225_mask = 1'h1;
  assign cache_v__T_225_en = reset;
  assign cache_v__T_226_data = 1'h0;
  assign cache_v__T_226_addr = 8'hd8;
  assign cache_v__T_226_mask = 1'h1;
  assign cache_v__T_226_en = reset;
  assign cache_v__T_227_data = 1'h0;
  assign cache_v__T_227_addr = 8'hd9;
  assign cache_v__T_227_mask = 1'h1;
  assign cache_v__T_227_en = reset;
  assign cache_v__T_228_data = 1'h0;
  assign cache_v__T_228_addr = 8'hda;
  assign cache_v__T_228_mask = 1'h1;
  assign cache_v__T_228_en = reset;
  assign cache_v__T_229_data = 1'h0;
  assign cache_v__T_229_addr = 8'hdb;
  assign cache_v__T_229_mask = 1'h1;
  assign cache_v__T_229_en = reset;
  assign cache_v__T_230_data = 1'h0;
  assign cache_v__T_230_addr = 8'hdc;
  assign cache_v__T_230_mask = 1'h1;
  assign cache_v__T_230_en = reset;
  assign cache_v__T_231_data = 1'h0;
  assign cache_v__T_231_addr = 8'hdd;
  assign cache_v__T_231_mask = 1'h1;
  assign cache_v__T_231_en = reset;
  assign cache_v__T_232_data = 1'h0;
  assign cache_v__T_232_addr = 8'hde;
  assign cache_v__T_232_mask = 1'h1;
  assign cache_v__T_232_en = reset;
  assign cache_v__T_233_data = 1'h0;
  assign cache_v__T_233_addr = 8'hdf;
  assign cache_v__T_233_mask = 1'h1;
  assign cache_v__T_233_en = reset;
  assign cache_v__T_234_data = 1'h0;
  assign cache_v__T_234_addr = 8'he0;
  assign cache_v__T_234_mask = 1'h1;
  assign cache_v__T_234_en = reset;
  assign cache_v__T_235_data = 1'h0;
  assign cache_v__T_235_addr = 8'he1;
  assign cache_v__T_235_mask = 1'h1;
  assign cache_v__T_235_en = reset;
  assign cache_v__T_236_data = 1'h0;
  assign cache_v__T_236_addr = 8'he2;
  assign cache_v__T_236_mask = 1'h1;
  assign cache_v__T_236_en = reset;
  assign cache_v__T_237_data = 1'h0;
  assign cache_v__T_237_addr = 8'he3;
  assign cache_v__T_237_mask = 1'h1;
  assign cache_v__T_237_en = reset;
  assign cache_v__T_238_data = 1'h0;
  assign cache_v__T_238_addr = 8'he4;
  assign cache_v__T_238_mask = 1'h1;
  assign cache_v__T_238_en = reset;
  assign cache_v__T_239_data = 1'h0;
  assign cache_v__T_239_addr = 8'he5;
  assign cache_v__T_239_mask = 1'h1;
  assign cache_v__T_239_en = reset;
  assign cache_v__T_240_data = 1'h0;
  assign cache_v__T_240_addr = 8'he6;
  assign cache_v__T_240_mask = 1'h1;
  assign cache_v__T_240_en = reset;
  assign cache_v__T_241_data = 1'h0;
  assign cache_v__T_241_addr = 8'he7;
  assign cache_v__T_241_mask = 1'h1;
  assign cache_v__T_241_en = reset;
  assign cache_v__T_242_data = 1'h0;
  assign cache_v__T_242_addr = 8'he8;
  assign cache_v__T_242_mask = 1'h1;
  assign cache_v__T_242_en = reset;
  assign cache_v__T_243_data = 1'h0;
  assign cache_v__T_243_addr = 8'he9;
  assign cache_v__T_243_mask = 1'h1;
  assign cache_v__T_243_en = reset;
  assign cache_v__T_244_data = 1'h0;
  assign cache_v__T_244_addr = 8'hea;
  assign cache_v__T_244_mask = 1'h1;
  assign cache_v__T_244_en = reset;
  assign cache_v__T_245_data = 1'h0;
  assign cache_v__T_245_addr = 8'heb;
  assign cache_v__T_245_mask = 1'h1;
  assign cache_v__T_245_en = reset;
  assign cache_v__T_246_data = 1'h0;
  assign cache_v__T_246_addr = 8'hec;
  assign cache_v__T_246_mask = 1'h1;
  assign cache_v__T_246_en = reset;
  assign cache_v__T_247_data = 1'h0;
  assign cache_v__T_247_addr = 8'hed;
  assign cache_v__T_247_mask = 1'h1;
  assign cache_v__T_247_en = reset;
  assign cache_v__T_248_data = 1'h0;
  assign cache_v__T_248_addr = 8'hee;
  assign cache_v__T_248_mask = 1'h1;
  assign cache_v__T_248_en = reset;
  assign cache_v__T_249_data = 1'h0;
  assign cache_v__T_249_addr = 8'hef;
  assign cache_v__T_249_mask = 1'h1;
  assign cache_v__T_249_en = reset;
  assign cache_v__T_250_data = 1'h0;
  assign cache_v__T_250_addr = 8'hf0;
  assign cache_v__T_250_mask = 1'h1;
  assign cache_v__T_250_en = reset;
  assign cache_v__T_251_data = 1'h0;
  assign cache_v__T_251_addr = 8'hf1;
  assign cache_v__T_251_mask = 1'h1;
  assign cache_v__T_251_en = reset;
  assign cache_v__T_252_data = 1'h0;
  assign cache_v__T_252_addr = 8'hf2;
  assign cache_v__T_252_mask = 1'h1;
  assign cache_v__T_252_en = reset;
  assign cache_v__T_253_data = 1'h0;
  assign cache_v__T_253_addr = 8'hf3;
  assign cache_v__T_253_mask = 1'h1;
  assign cache_v__T_253_en = reset;
  assign cache_v__T_254_data = 1'h0;
  assign cache_v__T_254_addr = 8'hf4;
  assign cache_v__T_254_mask = 1'h1;
  assign cache_v__T_254_en = reset;
  assign cache_v__T_255_data = 1'h0;
  assign cache_v__T_255_addr = 8'hf5;
  assign cache_v__T_255_mask = 1'h1;
  assign cache_v__T_255_en = reset;
  assign cache_v__T_256_data = 1'h0;
  assign cache_v__T_256_addr = 8'hf6;
  assign cache_v__T_256_mask = 1'h1;
  assign cache_v__T_256_en = reset;
  assign cache_v__T_257_data = 1'h0;
  assign cache_v__T_257_addr = 8'hf7;
  assign cache_v__T_257_mask = 1'h1;
  assign cache_v__T_257_en = reset;
  assign cache_v__T_258_data = 1'h0;
  assign cache_v__T_258_addr = 8'hf8;
  assign cache_v__T_258_mask = 1'h1;
  assign cache_v__T_258_en = reset;
  assign cache_v__T_259_data = 1'h0;
  assign cache_v__T_259_addr = 8'hf9;
  assign cache_v__T_259_mask = 1'h1;
  assign cache_v__T_259_en = reset;
  assign cache_v__T_260_data = 1'h0;
  assign cache_v__T_260_addr = 8'hfa;
  assign cache_v__T_260_mask = 1'h1;
  assign cache_v__T_260_en = reset;
  assign cache_v__T_261_data = 1'h0;
  assign cache_v__T_261_addr = 8'hfb;
  assign cache_v__T_261_mask = 1'h1;
  assign cache_v__T_261_en = reset;
  assign cache_v__T_262_data = 1'h0;
  assign cache_v__T_262_addr = 8'hfc;
  assign cache_v__T_262_mask = 1'h1;
  assign cache_v__T_262_en = reset;
  assign cache_v__T_263_data = 1'h0;
  assign cache_v__T_263_addr = 8'hfd;
  assign cache_v__T_263_mask = 1'h1;
  assign cache_v__T_263_en = reset;
  assign cache_v__T_264_data = 1'h0;
  assign cache_v__T_264_addr = 8'hfe;
  assign cache_v__T_264_mask = 1'h1;
  assign cache_v__T_264_en = reset;
  assign cache_v__T_265_data = 1'h0;
  assign cache_v__T_265_addr = 8'hff;
  assign cache_v__T_265_mask = 1'h1;
  assign cache_v__T_265_en = reset;
  assign cache_v_s1_entry_w_data = 1'h1;
  assign cache_v_s1_entry_w_addr = s1_in_addr[7:0];
  assign cache_v_s1_entry_w_mask = s1_resp & _T_285;
  assign cache_v_s1_entry_w_en = s1_resp & _T_285;
  assign cache_tag_s1_entry_r_addr = s1_in_addr[7:0];
  assign cache_tag_s1_entry_r_data = cache_tag[cache_tag_s1_entry_r_addr]; // @[icache.scala 91:18]
  assign cache_tag__T_8_data = 24'h0;
  assign cache_tag__T_8_addr = _T_6[7:0];
  assign cache_tag__T_8_mask = 1'h0;
  assign cache_tag__T_8_en = _T_1 & _T_5;
  assign cache_tag__T_10_data = 24'h0;
  assign cache_tag__T_10_addr = 8'h0;
  assign cache_tag__T_10_mask = 1'h0;
  assign cache_tag__T_10_en = reset;
  assign cache_tag__T_11_data = 24'h0;
  assign cache_tag__T_11_addr = 8'h1;
  assign cache_tag__T_11_mask = 1'h0;
  assign cache_tag__T_11_en = reset;
  assign cache_tag__T_12_data = 24'h0;
  assign cache_tag__T_12_addr = 8'h2;
  assign cache_tag__T_12_mask = 1'h0;
  assign cache_tag__T_12_en = reset;
  assign cache_tag__T_13_data = 24'h0;
  assign cache_tag__T_13_addr = 8'h3;
  assign cache_tag__T_13_mask = 1'h0;
  assign cache_tag__T_13_en = reset;
  assign cache_tag__T_14_data = 24'h0;
  assign cache_tag__T_14_addr = 8'h4;
  assign cache_tag__T_14_mask = 1'h0;
  assign cache_tag__T_14_en = reset;
  assign cache_tag__T_15_data = 24'h0;
  assign cache_tag__T_15_addr = 8'h5;
  assign cache_tag__T_15_mask = 1'h0;
  assign cache_tag__T_15_en = reset;
  assign cache_tag__T_16_data = 24'h0;
  assign cache_tag__T_16_addr = 8'h6;
  assign cache_tag__T_16_mask = 1'h0;
  assign cache_tag__T_16_en = reset;
  assign cache_tag__T_17_data = 24'h0;
  assign cache_tag__T_17_addr = 8'h7;
  assign cache_tag__T_17_mask = 1'h0;
  assign cache_tag__T_17_en = reset;
  assign cache_tag__T_18_data = 24'h0;
  assign cache_tag__T_18_addr = 8'h8;
  assign cache_tag__T_18_mask = 1'h0;
  assign cache_tag__T_18_en = reset;
  assign cache_tag__T_19_data = 24'h0;
  assign cache_tag__T_19_addr = 8'h9;
  assign cache_tag__T_19_mask = 1'h0;
  assign cache_tag__T_19_en = reset;
  assign cache_tag__T_20_data = 24'h0;
  assign cache_tag__T_20_addr = 8'ha;
  assign cache_tag__T_20_mask = 1'h0;
  assign cache_tag__T_20_en = reset;
  assign cache_tag__T_21_data = 24'h0;
  assign cache_tag__T_21_addr = 8'hb;
  assign cache_tag__T_21_mask = 1'h0;
  assign cache_tag__T_21_en = reset;
  assign cache_tag__T_22_data = 24'h0;
  assign cache_tag__T_22_addr = 8'hc;
  assign cache_tag__T_22_mask = 1'h0;
  assign cache_tag__T_22_en = reset;
  assign cache_tag__T_23_data = 24'h0;
  assign cache_tag__T_23_addr = 8'hd;
  assign cache_tag__T_23_mask = 1'h0;
  assign cache_tag__T_23_en = reset;
  assign cache_tag__T_24_data = 24'h0;
  assign cache_tag__T_24_addr = 8'he;
  assign cache_tag__T_24_mask = 1'h0;
  assign cache_tag__T_24_en = reset;
  assign cache_tag__T_25_data = 24'h0;
  assign cache_tag__T_25_addr = 8'hf;
  assign cache_tag__T_25_mask = 1'h0;
  assign cache_tag__T_25_en = reset;
  assign cache_tag__T_26_data = 24'h0;
  assign cache_tag__T_26_addr = 8'h10;
  assign cache_tag__T_26_mask = 1'h0;
  assign cache_tag__T_26_en = reset;
  assign cache_tag__T_27_data = 24'h0;
  assign cache_tag__T_27_addr = 8'h11;
  assign cache_tag__T_27_mask = 1'h0;
  assign cache_tag__T_27_en = reset;
  assign cache_tag__T_28_data = 24'h0;
  assign cache_tag__T_28_addr = 8'h12;
  assign cache_tag__T_28_mask = 1'h0;
  assign cache_tag__T_28_en = reset;
  assign cache_tag__T_29_data = 24'h0;
  assign cache_tag__T_29_addr = 8'h13;
  assign cache_tag__T_29_mask = 1'h0;
  assign cache_tag__T_29_en = reset;
  assign cache_tag__T_30_data = 24'h0;
  assign cache_tag__T_30_addr = 8'h14;
  assign cache_tag__T_30_mask = 1'h0;
  assign cache_tag__T_30_en = reset;
  assign cache_tag__T_31_data = 24'h0;
  assign cache_tag__T_31_addr = 8'h15;
  assign cache_tag__T_31_mask = 1'h0;
  assign cache_tag__T_31_en = reset;
  assign cache_tag__T_32_data = 24'h0;
  assign cache_tag__T_32_addr = 8'h16;
  assign cache_tag__T_32_mask = 1'h0;
  assign cache_tag__T_32_en = reset;
  assign cache_tag__T_33_data = 24'h0;
  assign cache_tag__T_33_addr = 8'h17;
  assign cache_tag__T_33_mask = 1'h0;
  assign cache_tag__T_33_en = reset;
  assign cache_tag__T_34_data = 24'h0;
  assign cache_tag__T_34_addr = 8'h18;
  assign cache_tag__T_34_mask = 1'h0;
  assign cache_tag__T_34_en = reset;
  assign cache_tag__T_35_data = 24'h0;
  assign cache_tag__T_35_addr = 8'h19;
  assign cache_tag__T_35_mask = 1'h0;
  assign cache_tag__T_35_en = reset;
  assign cache_tag__T_36_data = 24'h0;
  assign cache_tag__T_36_addr = 8'h1a;
  assign cache_tag__T_36_mask = 1'h0;
  assign cache_tag__T_36_en = reset;
  assign cache_tag__T_37_data = 24'h0;
  assign cache_tag__T_37_addr = 8'h1b;
  assign cache_tag__T_37_mask = 1'h0;
  assign cache_tag__T_37_en = reset;
  assign cache_tag__T_38_data = 24'h0;
  assign cache_tag__T_38_addr = 8'h1c;
  assign cache_tag__T_38_mask = 1'h0;
  assign cache_tag__T_38_en = reset;
  assign cache_tag__T_39_data = 24'h0;
  assign cache_tag__T_39_addr = 8'h1d;
  assign cache_tag__T_39_mask = 1'h0;
  assign cache_tag__T_39_en = reset;
  assign cache_tag__T_40_data = 24'h0;
  assign cache_tag__T_40_addr = 8'h1e;
  assign cache_tag__T_40_mask = 1'h0;
  assign cache_tag__T_40_en = reset;
  assign cache_tag__T_41_data = 24'h0;
  assign cache_tag__T_41_addr = 8'h1f;
  assign cache_tag__T_41_mask = 1'h0;
  assign cache_tag__T_41_en = reset;
  assign cache_tag__T_42_data = 24'h0;
  assign cache_tag__T_42_addr = 8'h20;
  assign cache_tag__T_42_mask = 1'h0;
  assign cache_tag__T_42_en = reset;
  assign cache_tag__T_43_data = 24'h0;
  assign cache_tag__T_43_addr = 8'h21;
  assign cache_tag__T_43_mask = 1'h0;
  assign cache_tag__T_43_en = reset;
  assign cache_tag__T_44_data = 24'h0;
  assign cache_tag__T_44_addr = 8'h22;
  assign cache_tag__T_44_mask = 1'h0;
  assign cache_tag__T_44_en = reset;
  assign cache_tag__T_45_data = 24'h0;
  assign cache_tag__T_45_addr = 8'h23;
  assign cache_tag__T_45_mask = 1'h0;
  assign cache_tag__T_45_en = reset;
  assign cache_tag__T_46_data = 24'h0;
  assign cache_tag__T_46_addr = 8'h24;
  assign cache_tag__T_46_mask = 1'h0;
  assign cache_tag__T_46_en = reset;
  assign cache_tag__T_47_data = 24'h0;
  assign cache_tag__T_47_addr = 8'h25;
  assign cache_tag__T_47_mask = 1'h0;
  assign cache_tag__T_47_en = reset;
  assign cache_tag__T_48_data = 24'h0;
  assign cache_tag__T_48_addr = 8'h26;
  assign cache_tag__T_48_mask = 1'h0;
  assign cache_tag__T_48_en = reset;
  assign cache_tag__T_49_data = 24'h0;
  assign cache_tag__T_49_addr = 8'h27;
  assign cache_tag__T_49_mask = 1'h0;
  assign cache_tag__T_49_en = reset;
  assign cache_tag__T_50_data = 24'h0;
  assign cache_tag__T_50_addr = 8'h28;
  assign cache_tag__T_50_mask = 1'h0;
  assign cache_tag__T_50_en = reset;
  assign cache_tag__T_51_data = 24'h0;
  assign cache_tag__T_51_addr = 8'h29;
  assign cache_tag__T_51_mask = 1'h0;
  assign cache_tag__T_51_en = reset;
  assign cache_tag__T_52_data = 24'h0;
  assign cache_tag__T_52_addr = 8'h2a;
  assign cache_tag__T_52_mask = 1'h0;
  assign cache_tag__T_52_en = reset;
  assign cache_tag__T_53_data = 24'h0;
  assign cache_tag__T_53_addr = 8'h2b;
  assign cache_tag__T_53_mask = 1'h0;
  assign cache_tag__T_53_en = reset;
  assign cache_tag__T_54_data = 24'h0;
  assign cache_tag__T_54_addr = 8'h2c;
  assign cache_tag__T_54_mask = 1'h0;
  assign cache_tag__T_54_en = reset;
  assign cache_tag__T_55_data = 24'h0;
  assign cache_tag__T_55_addr = 8'h2d;
  assign cache_tag__T_55_mask = 1'h0;
  assign cache_tag__T_55_en = reset;
  assign cache_tag__T_56_data = 24'h0;
  assign cache_tag__T_56_addr = 8'h2e;
  assign cache_tag__T_56_mask = 1'h0;
  assign cache_tag__T_56_en = reset;
  assign cache_tag__T_57_data = 24'h0;
  assign cache_tag__T_57_addr = 8'h2f;
  assign cache_tag__T_57_mask = 1'h0;
  assign cache_tag__T_57_en = reset;
  assign cache_tag__T_58_data = 24'h0;
  assign cache_tag__T_58_addr = 8'h30;
  assign cache_tag__T_58_mask = 1'h0;
  assign cache_tag__T_58_en = reset;
  assign cache_tag__T_59_data = 24'h0;
  assign cache_tag__T_59_addr = 8'h31;
  assign cache_tag__T_59_mask = 1'h0;
  assign cache_tag__T_59_en = reset;
  assign cache_tag__T_60_data = 24'h0;
  assign cache_tag__T_60_addr = 8'h32;
  assign cache_tag__T_60_mask = 1'h0;
  assign cache_tag__T_60_en = reset;
  assign cache_tag__T_61_data = 24'h0;
  assign cache_tag__T_61_addr = 8'h33;
  assign cache_tag__T_61_mask = 1'h0;
  assign cache_tag__T_61_en = reset;
  assign cache_tag__T_62_data = 24'h0;
  assign cache_tag__T_62_addr = 8'h34;
  assign cache_tag__T_62_mask = 1'h0;
  assign cache_tag__T_62_en = reset;
  assign cache_tag__T_63_data = 24'h0;
  assign cache_tag__T_63_addr = 8'h35;
  assign cache_tag__T_63_mask = 1'h0;
  assign cache_tag__T_63_en = reset;
  assign cache_tag__T_64_data = 24'h0;
  assign cache_tag__T_64_addr = 8'h36;
  assign cache_tag__T_64_mask = 1'h0;
  assign cache_tag__T_64_en = reset;
  assign cache_tag__T_65_data = 24'h0;
  assign cache_tag__T_65_addr = 8'h37;
  assign cache_tag__T_65_mask = 1'h0;
  assign cache_tag__T_65_en = reset;
  assign cache_tag__T_66_data = 24'h0;
  assign cache_tag__T_66_addr = 8'h38;
  assign cache_tag__T_66_mask = 1'h0;
  assign cache_tag__T_66_en = reset;
  assign cache_tag__T_67_data = 24'h0;
  assign cache_tag__T_67_addr = 8'h39;
  assign cache_tag__T_67_mask = 1'h0;
  assign cache_tag__T_67_en = reset;
  assign cache_tag__T_68_data = 24'h0;
  assign cache_tag__T_68_addr = 8'h3a;
  assign cache_tag__T_68_mask = 1'h0;
  assign cache_tag__T_68_en = reset;
  assign cache_tag__T_69_data = 24'h0;
  assign cache_tag__T_69_addr = 8'h3b;
  assign cache_tag__T_69_mask = 1'h0;
  assign cache_tag__T_69_en = reset;
  assign cache_tag__T_70_data = 24'h0;
  assign cache_tag__T_70_addr = 8'h3c;
  assign cache_tag__T_70_mask = 1'h0;
  assign cache_tag__T_70_en = reset;
  assign cache_tag__T_71_data = 24'h0;
  assign cache_tag__T_71_addr = 8'h3d;
  assign cache_tag__T_71_mask = 1'h0;
  assign cache_tag__T_71_en = reset;
  assign cache_tag__T_72_data = 24'h0;
  assign cache_tag__T_72_addr = 8'h3e;
  assign cache_tag__T_72_mask = 1'h0;
  assign cache_tag__T_72_en = reset;
  assign cache_tag__T_73_data = 24'h0;
  assign cache_tag__T_73_addr = 8'h3f;
  assign cache_tag__T_73_mask = 1'h0;
  assign cache_tag__T_73_en = reset;
  assign cache_tag__T_74_data = 24'h0;
  assign cache_tag__T_74_addr = 8'h40;
  assign cache_tag__T_74_mask = 1'h0;
  assign cache_tag__T_74_en = reset;
  assign cache_tag__T_75_data = 24'h0;
  assign cache_tag__T_75_addr = 8'h41;
  assign cache_tag__T_75_mask = 1'h0;
  assign cache_tag__T_75_en = reset;
  assign cache_tag__T_76_data = 24'h0;
  assign cache_tag__T_76_addr = 8'h42;
  assign cache_tag__T_76_mask = 1'h0;
  assign cache_tag__T_76_en = reset;
  assign cache_tag__T_77_data = 24'h0;
  assign cache_tag__T_77_addr = 8'h43;
  assign cache_tag__T_77_mask = 1'h0;
  assign cache_tag__T_77_en = reset;
  assign cache_tag__T_78_data = 24'h0;
  assign cache_tag__T_78_addr = 8'h44;
  assign cache_tag__T_78_mask = 1'h0;
  assign cache_tag__T_78_en = reset;
  assign cache_tag__T_79_data = 24'h0;
  assign cache_tag__T_79_addr = 8'h45;
  assign cache_tag__T_79_mask = 1'h0;
  assign cache_tag__T_79_en = reset;
  assign cache_tag__T_80_data = 24'h0;
  assign cache_tag__T_80_addr = 8'h46;
  assign cache_tag__T_80_mask = 1'h0;
  assign cache_tag__T_80_en = reset;
  assign cache_tag__T_81_data = 24'h0;
  assign cache_tag__T_81_addr = 8'h47;
  assign cache_tag__T_81_mask = 1'h0;
  assign cache_tag__T_81_en = reset;
  assign cache_tag__T_82_data = 24'h0;
  assign cache_tag__T_82_addr = 8'h48;
  assign cache_tag__T_82_mask = 1'h0;
  assign cache_tag__T_82_en = reset;
  assign cache_tag__T_83_data = 24'h0;
  assign cache_tag__T_83_addr = 8'h49;
  assign cache_tag__T_83_mask = 1'h0;
  assign cache_tag__T_83_en = reset;
  assign cache_tag__T_84_data = 24'h0;
  assign cache_tag__T_84_addr = 8'h4a;
  assign cache_tag__T_84_mask = 1'h0;
  assign cache_tag__T_84_en = reset;
  assign cache_tag__T_85_data = 24'h0;
  assign cache_tag__T_85_addr = 8'h4b;
  assign cache_tag__T_85_mask = 1'h0;
  assign cache_tag__T_85_en = reset;
  assign cache_tag__T_86_data = 24'h0;
  assign cache_tag__T_86_addr = 8'h4c;
  assign cache_tag__T_86_mask = 1'h0;
  assign cache_tag__T_86_en = reset;
  assign cache_tag__T_87_data = 24'h0;
  assign cache_tag__T_87_addr = 8'h4d;
  assign cache_tag__T_87_mask = 1'h0;
  assign cache_tag__T_87_en = reset;
  assign cache_tag__T_88_data = 24'h0;
  assign cache_tag__T_88_addr = 8'h4e;
  assign cache_tag__T_88_mask = 1'h0;
  assign cache_tag__T_88_en = reset;
  assign cache_tag__T_89_data = 24'h0;
  assign cache_tag__T_89_addr = 8'h4f;
  assign cache_tag__T_89_mask = 1'h0;
  assign cache_tag__T_89_en = reset;
  assign cache_tag__T_90_data = 24'h0;
  assign cache_tag__T_90_addr = 8'h50;
  assign cache_tag__T_90_mask = 1'h0;
  assign cache_tag__T_90_en = reset;
  assign cache_tag__T_91_data = 24'h0;
  assign cache_tag__T_91_addr = 8'h51;
  assign cache_tag__T_91_mask = 1'h0;
  assign cache_tag__T_91_en = reset;
  assign cache_tag__T_92_data = 24'h0;
  assign cache_tag__T_92_addr = 8'h52;
  assign cache_tag__T_92_mask = 1'h0;
  assign cache_tag__T_92_en = reset;
  assign cache_tag__T_93_data = 24'h0;
  assign cache_tag__T_93_addr = 8'h53;
  assign cache_tag__T_93_mask = 1'h0;
  assign cache_tag__T_93_en = reset;
  assign cache_tag__T_94_data = 24'h0;
  assign cache_tag__T_94_addr = 8'h54;
  assign cache_tag__T_94_mask = 1'h0;
  assign cache_tag__T_94_en = reset;
  assign cache_tag__T_95_data = 24'h0;
  assign cache_tag__T_95_addr = 8'h55;
  assign cache_tag__T_95_mask = 1'h0;
  assign cache_tag__T_95_en = reset;
  assign cache_tag__T_96_data = 24'h0;
  assign cache_tag__T_96_addr = 8'h56;
  assign cache_tag__T_96_mask = 1'h0;
  assign cache_tag__T_96_en = reset;
  assign cache_tag__T_97_data = 24'h0;
  assign cache_tag__T_97_addr = 8'h57;
  assign cache_tag__T_97_mask = 1'h0;
  assign cache_tag__T_97_en = reset;
  assign cache_tag__T_98_data = 24'h0;
  assign cache_tag__T_98_addr = 8'h58;
  assign cache_tag__T_98_mask = 1'h0;
  assign cache_tag__T_98_en = reset;
  assign cache_tag__T_99_data = 24'h0;
  assign cache_tag__T_99_addr = 8'h59;
  assign cache_tag__T_99_mask = 1'h0;
  assign cache_tag__T_99_en = reset;
  assign cache_tag__T_100_data = 24'h0;
  assign cache_tag__T_100_addr = 8'h5a;
  assign cache_tag__T_100_mask = 1'h0;
  assign cache_tag__T_100_en = reset;
  assign cache_tag__T_101_data = 24'h0;
  assign cache_tag__T_101_addr = 8'h5b;
  assign cache_tag__T_101_mask = 1'h0;
  assign cache_tag__T_101_en = reset;
  assign cache_tag__T_102_data = 24'h0;
  assign cache_tag__T_102_addr = 8'h5c;
  assign cache_tag__T_102_mask = 1'h0;
  assign cache_tag__T_102_en = reset;
  assign cache_tag__T_103_data = 24'h0;
  assign cache_tag__T_103_addr = 8'h5d;
  assign cache_tag__T_103_mask = 1'h0;
  assign cache_tag__T_103_en = reset;
  assign cache_tag__T_104_data = 24'h0;
  assign cache_tag__T_104_addr = 8'h5e;
  assign cache_tag__T_104_mask = 1'h0;
  assign cache_tag__T_104_en = reset;
  assign cache_tag__T_105_data = 24'h0;
  assign cache_tag__T_105_addr = 8'h5f;
  assign cache_tag__T_105_mask = 1'h0;
  assign cache_tag__T_105_en = reset;
  assign cache_tag__T_106_data = 24'h0;
  assign cache_tag__T_106_addr = 8'h60;
  assign cache_tag__T_106_mask = 1'h0;
  assign cache_tag__T_106_en = reset;
  assign cache_tag__T_107_data = 24'h0;
  assign cache_tag__T_107_addr = 8'h61;
  assign cache_tag__T_107_mask = 1'h0;
  assign cache_tag__T_107_en = reset;
  assign cache_tag__T_108_data = 24'h0;
  assign cache_tag__T_108_addr = 8'h62;
  assign cache_tag__T_108_mask = 1'h0;
  assign cache_tag__T_108_en = reset;
  assign cache_tag__T_109_data = 24'h0;
  assign cache_tag__T_109_addr = 8'h63;
  assign cache_tag__T_109_mask = 1'h0;
  assign cache_tag__T_109_en = reset;
  assign cache_tag__T_110_data = 24'h0;
  assign cache_tag__T_110_addr = 8'h64;
  assign cache_tag__T_110_mask = 1'h0;
  assign cache_tag__T_110_en = reset;
  assign cache_tag__T_111_data = 24'h0;
  assign cache_tag__T_111_addr = 8'h65;
  assign cache_tag__T_111_mask = 1'h0;
  assign cache_tag__T_111_en = reset;
  assign cache_tag__T_112_data = 24'h0;
  assign cache_tag__T_112_addr = 8'h66;
  assign cache_tag__T_112_mask = 1'h0;
  assign cache_tag__T_112_en = reset;
  assign cache_tag__T_113_data = 24'h0;
  assign cache_tag__T_113_addr = 8'h67;
  assign cache_tag__T_113_mask = 1'h0;
  assign cache_tag__T_113_en = reset;
  assign cache_tag__T_114_data = 24'h0;
  assign cache_tag__T_114_addr = 8'h68;
  assign cache_tag__T_114_mask = 1'h0;
  assign cache_tag__T_114_en = reset;
  assign cache_tag__T_115_data = 24'h0;
  assign cache_tag__T_115_addr = 8'h69;
  assign cache_tag__T_115_mask = 1'h0;
  assign cache_tag__T_115_en = reset;
  assign cache_tag__T_116_data = 24'h0;
  assign cache_tag__T_116_addr = 8'h6a;
  assign cache_tag__T_116_mask = 1'h0;
  assign cache_tag__T_116_en = reset;
  assign cache_tag__T_117_data = 24'h0;
  assign cache_tag__T_117_addr = 8'h6b;
  assign cache_tag__T_117_mask = 1'h0;
  assign cache_tag__T_117_en = reset;
  assign cache_tag__T_118_data = 24'h0;
  assign cache_tag__T_118_addr = 8'h6c;
  assign cache_tag__T_118_mask = 1'h0;
  assign cache_tag__T_118_en = reset;
  assign cache_tag__T_119_data = 24'h0;
  assign cache_tag__T_119_addr = 8'h6d;
  assign cache_tag__T_119_mask = 1'h0;
  assign cache_tag__T_119_en = reset;
  assign cache_tag__T_120_data = 24'h0;
  assign cache_tag__T_120_addr = 8'h6e;
  assign cache_tag__T_120_mask = 1'h0;
  assign cache_tag__T_120_en = reset;
  assign cache_tag__T_121_data = 24'h0;
  assign cache_tag__T_121_addr = 8'h6f;
  assign cache_tag__T_121_mask = 1'h0;
  assign cache_tag__T_121_en = reset;
  assign cache_tag__T_122_data = 24'h0;
  assign cache_tag__T_122_addr = 8'h70;
  assign cache_tag__T_122_mask = 1'h0;
  assign cache_tag__T_122_en = reset;
  assign cache_tag__T_123_data = 24'h0;
  assign cache_tag__T_123_addr = 8'h71;
  assign cache_tag__T_123_mask = 1'h0;
  assign cache_tag__T_123_en = reset;
  assign cache_tag__T_124_data = 24'h0;
  assign cache_tag__T_124_addr = 8'h72;
  assign cache_tag__T_124_mask = 1'h0;
  assign cache_tag__T_124_en = reset;
  assign cache_tag__T_125_data = 24'h0;
  assign cache_tag__T_125_addr = 8'h73;
  assign cache_tag__T_125_mask = 1'h0;
  assign cache_tag__T_125_en = reset;
  assign cache_tag__T_126_data = 24'h0;
  assign cache_tag__T_126_addr = 8'h74;
  assign cache_tag__T_126_mask = 1'h0;
  assign cache_tag__T_126_en = reset;
  assign cache_tag__T_127_data = 24'h0;
  assign cache_tag__T_127_addr = 8'h75;
  assign cache_tag__T_127_mask = 1'h0;
  assign cache_tag__T_127_en = reset;
  assign cache_tag__T_128_data = 24'h0;
  assign cache_tag__T_128_addr = 8'h76;
  assign cache_tag__T_128_mask = 1'h0;
  assign cache_tag__T_128_en = reset;
  assign cache_tag__T_129_data = 24'h0;
  assign cache_tag__T_129_addr = 8'h77;
  assign cache_tag__T_129_mask = 1'h0;
  assign cache_tag__T_129_en = reset;
  assign cache_tag__T_130_data = 24'h0;
  assign cache_tag__T_130_addr = 8'h78;
  assign cache_tag__T_130_mask = 1'h0;
  assign cache_tag__T_130_en = reset;
  assign cache_tag__T_131_data = 24'h0;
  assign cache_tag__T_131_addr = 8'h79;
  assign cache_tag__T_131_mask = 1'h0;
  assign cache_tag__T_131_en = reset;
  assign cache_tag__T_132_data = 24'h0;
  assign cache_tag__T_132_addr = 8'h7a;
  assign cache_tag__T_132_mask = 1'h0;
  assign cache_tag__T_132_en = reset;
  assign cache_tag__T_133_data = 24'h0;
  assign cache_tag__T_133_addr = 8'h7b;
  assign cache_tag__T_133_mask = 1'h0;
  assign cache_tag__T_133_en = reset;
  assign cache_tag__T_134_data = 24'h0;
  assign cache_tag__T_134_addr = 8'h7c;
  assign cache_tag__T_134_mask = 1'h0;
  assign cache_tag__T_134_en = reset;
  assign cache_tag__T_135_data = 24'h0;
  assign cache_tag__T_135_addr = 8'h7d;
  assign cache_tag__T_135_mask = 1'h0;
  assign cache_tag__T_135_en = reset;
  assign cache_tag__T_136_data = 24'h0;
  assign cache_tag__T_136_addr = 8'h7e;
  assign cache_tag__T_136_mask = 1'h0;
  assign cache_tag__T_136_en = reset;
  assign cache_tag__T_137_data = 24'h0;
  assign cache_tag__T_137_addr = 8'h7f;
  assign cache_tag__T_137_mask = 1'h0;
  assign cache_tag__T_137_en = reset;
  assign cache_tag__T_138_data = 24'h0;
  assign cache_tag__T_138_addr = 8'h80;
  assign cache_tag__T_138_mask = 1'h0;
  assign cache_tag__T_138_en = reset;
  assign cache_tag__T_139_data = 24'h0;
  assign cache_tag__T_139_addr = 8'h81;
  assign cache_tag__T_139_mask = 1'h0;
  assign cache_tag__T_139_en = reset;
  assign cache_tag__T_140_data = 24'h0;
  assign cache_tag__T_140_addr = 8'h82;
  assign cache_tag__T_140_mask = 1'h0;
  assign cache_tag__T_140_en = reset;
  assign cache_tag__T_141_data = 24'h0;
  assign cache_tag__T_141_addr = 8'h83;
  assign cache_tag__T_141_mask = 1'h0;
  assign cache_tag__T_141_en = reset;
  assign cache_tag__T_142_data = 24'h0;
  assign cache_tag__T_142_addr = 8'h84;
  assign cache_tag__T_142_mask = 1'h0;
  assign cache_tag__T_142_en = reset;
  assign cache_tag__T_143_data = 24'h0;
  assign cache_tag__T_143_addr = 8'h85;
  assign cache_tag__T_143_mask = 1'h0;
  assign cache_tag__T_143_en = reset;
  assign cache_tag__T_144_data = 24'h0;
  assign cache_tag__T_144_addr = 8'h86;
  assign cache_tag__T_144_mask = 1'h0;
  assign cache_tag__T_144_en = reset;
  assign cache_tag__T_145_data = 24'h0;
  assign cache_tag__T_145_addr = 8'h87;
  assign cache_tag__T_145_mask = 1'h0;
  assign cache_tag__T_145_en = reset;
  assign cache_tag__T_146_data = 24'h0;
  assign cache_tag__T_146_addr = 8'h88;
  assign cache_tag__T_146_mask = 1'h0;
  assign cache_tag__T_146_en = reset;
  assign cache_tag__T_147_data = 24'h0;
  assign cache_tag__T_147_addr = 8'h89;
  assign cache_tag__T_147_mask = 1'h0;
  assign cache_tag__T_147_en = reset;
  assign cache_tag__T_148_data = 24'h0;
  assign cache_tag__T_148_addr = 8'h8a;
  assign cache_tag__T_148_mask = 1'h0;
  assign cache_tag__T_148_en = reset;
  assign cache_tag__T_149_data = 24'h0;
  assign cache_tag__T_149_addr = 8'h8b;
  assign cache_tag__T_149_mask = 1'h0;
  assign cache_tag__T_149_en = reset;
  assign cache_tag__T_150_data = 24'h0;
  assign cache_tag__T_150_addr = 8'h8c;
  assign cache_tag__T_150_mask = 1'h0;
  assign cache_tag__T_150_en = reset;
  assign cache_tag__T_151_data = 24'h0;
  assign cache_tag__T_151_addr = 8'h8d;
  assign cache_tag__T_151_mask = 1'h0;
  assign cache_tag__T_151_en = reset;
  assign cache_tag__T_152_data = 24'h0;
  assign cache_tag__T_152_addr = 8'h8e;
  assign cache_tag__T_152_mask = 1'h0;
  assign cache_tag__T_152_en = reset;
  assign cache_tag__T_153_data = 24'h0;
  assign cache_tag__T_153_addr = 8'h8f;
  assign cache_tag__T_153_mask = 1'h0;
  assign cache_tag__T_153_en = reset;
  assign cache_tag__T_154_data = 24'h0;
  assign cache_tag__T_154_addr = 8'h90;
  assign cache_tag__T_154_mask = 1'h0;
  assign cache_tag__T_154_en = reset;
  assign cache_tag__T_155_data = 24'h0;
  assign cache_tag__T_155_addr = 8'h91;
  assign cache_tag__T_155_mask = 1'h0;
  assign cache_tag__T_155_en = reset;
  assign cache_tag__T_156_data = 24'h0;
  assign cache_tag__T_156_addr = 8'h92;
  assign cache_tag__T_156_mask = 1'h0;
  assign cache_tag__T_156_en = reset;
  assign cache_tag__T_157_data = 24'h0;
  assign cache_tag__T_157_addr = 8'h93;
  assign cache_tag__T_157_mask = 1'h0;
  assign cache_tag__T_157_en = reset;
  assign cache_tag__T_158_data = 24'h0;
  assign cache_tag__T_158_addr = 8'h94;
  assign cache_tag__T_158_mask = 1'h0;
  assign cache_tag__T_158_en = reset;
  assign cache_tag__T_159_data = 24'h0;
  assign cache_tag__T_159_addr = 8'h95;
  assign cache_tag__T_159_mask = 1'h0;
  assign cache_tag__T_159_en = reset;
  assign cache_tag__T_160_data = 24'h0;
  assign cache_tag__T_160_addr = 8'h96;
  assign cache_tag__T_160_mask = 1'h0;
  assign cache_tag__T_160_en = reset;
  assign cache_tag__T_161_data = 24'h0;
  assign cache_tag__T_161_addr = 8'h97;
  assign cache_tag__T_161_mask = 1'h0;
  assign cache_tag__T_161_en = reset;
  assign cache_tag__T_162_data = 24'h0;
  assign cache_tag__T_162_addr = 8'h98;
  assign cache_tag__T_162_mask = 1'h0;
  assign cache_tag__T_162_en = reset;
  assign cache_tag__T_163_data = 24'h0;
  assign cache_tag__T_163_addr = 8'h99;
  assign cache_tag__T_163_mask = 1'h0;
  assign cache_tag__T_163_en = reset;
  assign cache_tag__T_164_data = 24'h0;
  assign cache_tag__T_164_addr = 8'h9a;
  assign cache_tag__T_164_mask = 1'h0;
  assign cache_tag__T_164_en = reset;
  assign cache_tag__T_165_data = 24'h0;
  assign cache_tag__T_165_addr = 8'h9b;
  assign cache_tag__T_165_mask = 1'h0;
  assign cache_tag__T_165_en = reset;
  assign cache_tag__T_166_data = 24'h0;
  assign cache_tag__T_166_addr = 8'h9c;
  assign cache_tag__T_166_mask = 1'h0;
  assign cache_tag__T_166_en = reset;
  assign cache_tag__T_167_data = 24'h0;
  assign cache_tag__T_167_addr = 8'h9d;
  assign cache_tag__T_167_mask = 1'h0;
  assign cache_tag__T_167_en = reset;
  assign cache_tag__T_168_data = 24'h0;
  assign cache_tag__T_168_addr = 8'h9e;
  assign cache_tag__T_168_mask = 1'h0;
  assign cache_tag__T_168_en = reset;
  assign cache_tag__T_169_data = 24'h0;
  assign cache_tag__T_169_addr = 8'h9f;
  assign cache_tag__T_169_mask = 1'h0;
  assign cache_tag__T_169_en = reset;
  assign cache_tag__T_170_data = 24'h0;
  assign cache_tag__T_170_addr = 8'ha0;
  assign cache_tag__T_170_mask = 1'h0;
  assign cache_tag__T_170_en = reset;
  assign cache_tag__T_171_data = 24'h0;
  assign cache_tag__T_171_addr = 8'ha1;
  assign cache_tag__T_171_mask = 1'h0;
  assign cache_tag__T_171_en = reset;
  assign cache_tag__T_172_data = 24'h0;
  assign cache_tag__T_172_addr = 8'ha2;
  assign cache_tag__T_172_mask = 1'h0;
  assign cache_tag__T_172_en = reset;
  assign cache_tag__T_173_data = 24'h0;
  assign cache_tag__T_173_addr = 8'ha3;
  assign cache_tag__T_173_mask = 1'h0;
  assign cache_tag__T_173_en = reset;
  assign cache_tag__T_174_data = 24'h0;
  assign cache_tag__T_174_addr = 8'ha4;
  assign cache_tag__T_174_mask = 1'h0;
  assign cache_tag__T_174_en = reset;
  assign cache_tag__T_175_data = 24'h0;
  assign cache_tag__T_175_addr = 8'ha5;
  assign cache_tag__T_175_mask = 1'h0;
  assign cache_tag__T_175_en = reset;
  assign cache_tag__T_176_data = 24'h0;
  assign cache_tag__T_176_addr = 8'ha6;
  assign cache_tag__T_176_mask = 1'h0;
  assign cache_tag__T_176_en = reset;
  assign cache_tag__T_177_data = 24'h0;
  assign cache_tag__T_177_addr = 8'ha7;
  assign cache_tag__T_177_mask = 1'h0;
  assign cache_tag__T_177_en = reset;
  assign cache_tag__T_178_data = 24'h0;
  assign cache_tag__T_178_addr = 8'ha8;
  assign cache_tag__T_178_mask = 1'h0;
  assign cache_tag__T_178_en = reset;
  assign cache_tag__T_179_data = 24'h0;
  assign cache_tag__T_179_addr = 8'ha9;
  assign cache_tag__T_179_mask = 1'h0;
  assign cache_tag__T_179_en = reset;
  assign cache_tag__T_180_data = 24'h0;
  assign cache_tag__T_180_addr = 8'haa;
  assign cache_tag__T_180_mask = 1'h0;
  assign cache_tag__T_180_en = reset;
  assign cache_tag__T_181_data = 24'h0;
  assign cache_tag__T_181_addr = 8'hab;
  assign cache_tag__T_181_mask = 1'h0;
  assign cache_tag__T_181_en = reset;
  assign cache_tag__T_182_data = 24'h0;
  assign cache_tag__T_182_addr = 8'hac;
  assign cache_tag__T_182_mask = 1'h0;
  assign cache_tag__T_182_en = reset;
  assign cache_tag__T_183_data = 24'h0;
  assign cache_tag__T_183_addr = 8'had;
  assign cache_tag__T_183_mask = 1'h0;
  assign cache_tag__T_183_en = reset;
  assign cache_tag__T_184_data = 24'h0;
  assign cache_tag__T_184_addr = 8'hae;
  assign cache_tag__T_184_mask = 1'h0;
  assign cache_tag__T_184_en = reset;
  assign cache_tag__T_185_data = 24'h0;
  assign cache_tag__T_185_addr = 8'haf;
  assign cache_tag__T_185_mask = 1'h0;
  assign cache_tag__T_185_en = reset;
  assign cache_tag__T_186_data = 24'h0;
  assign cache_tag__T_186_addr = 8'hb0;
  assign cache_tag__T_186_mask = 1'h0;
  assign cache_tag__T_186_en = reset;
  assign cache_tag__T_187_data = 24'h0;
  assign cache_tag__T_187_addr = 8'hb1;
  assign cache_tag__T_187_mask = 1'h0;
  assign cache_tag__T_187_en = reset;
  assign cache_tag__T_188_data = 24'h0;
  assign cache_tag__T_188_addr = 8'hb2;
  assign cache_tag__T_188_mask = 1'h0;
  assign cache_tag__T_188_en = reset;
  assign cache_tag__T_189_data = 24'h0;
  assign cache_tag__T_189_addr = 8'hb3;
  assign cache_tag__T_189_mask = 1'h0;
  assign cache_tag__T_189_en = reset;
  assign cache_tag__T_190_data = 24'h0;
  assign cache_tag__T_190_addr = 8'hb4;
  assign cache_tag__T_190_mask = 1'h0;
  assign cache_tag__T_190_en = reset;
  assign cache_tag__T_191_data = 24'h0;
  assign cache_tag__T_191_addr = 8'hb5;
  assign cache_tag__T_191_mask = 1'h0;
  assign cache_tag__T_191_en = reset;
  assign cache_tag__T_192_data = 24'h0;
  assign cache_tag__T_192_addr = 8'hb6;
  assign cache_tag__T_192_mask = 1'h0;
  assign cache_tag__T_192_en = reset;
  assign cache_tag__T_193_data = 24'h0;
  assign cache_tag__T_193_addr = 8'hb7;
  assign cache_tag__T_193_mask = 1'h0;
  assign cache_tag__T_193_en = reset;
  assign cache_tag__T_194_data = 24'h0;
  assign cache_tag__T_194_addr = 8'hb8;
  assign cache_tag__T_194_mask = 1'h0;
  assign cache_tag__T_194_en = reset;
  assign cache_tag__T_195_data = 24'h0;
  assign cache_tag__T_195_addr = 8'hb9;
  assign cache_tag__T_195_mask = 1'h0;
  assign cache_tag__T_195_en = reset;
  assign cache_tag__T_196_data = 24'h0;
  assign cache_tag__T_196_addr = 8'hba;
  assign cache_tag__T_196_mask = 1'h0;
  assign cache_tag__T_196_en = reset;
  assign cache_tag__T_197_data = 24'h0;
  assign cache_tag__T_197_addr = 8'hbb;
  assign cache_tag__T_197_mask = 1'h0;
  assign cache_tag__T_197_en = reset;
  assign cache_tag__T_198_data = 24'h0;
  assign cache_tag__T_198_addr = 8'hbc;
  assign cache_tag__T_198_mask = 1'h0;
  assign cache_tag__T_198_en = reset;
  assign cache_tag__T_199_data = 24'h0;
  assign cache_tag__T_199_addr = 8'hbd;
  assign cache_tag__T_199_mask = 1'h0;
  assign cache_tag__T_199_en = reset;
  assign cache_tag__T_200_data = 24'h0;
  assign cache_tag__T_200_addr = 8'hbe;
  assign cache_tag__T_200_mask = 1'h0;
  assign cache_tag__T_200_en = reset;
  assign cache_tag__T_201_data = 24'h0;
  assign cache_tag__T_201_addr = 8'hbf;
  assign cache_tag__T_201_mask = 1'h0;
  assign cache_tag__T_201_en = reset;
  assign cache_tag__T_202_data = 24'h0;
  assign cache_tag__T_202_addr = 8'hc0;
  assign cache_tag__T_202_mask = 1'h0;
  assign cache_tag__T_202_en = reset;
  assign cache_tag__T_203_data = 24'h0;
  assign cache_tag__T_203_addr = 8'hc1;
  assign cache_tag__T_203_mask = 1'h0;
  assign cache_tag__T_203_en = reset;
  assign cache_tag__T_204_data = 24'h0;
  assign cache_tag__T_204_addr = 8'hc2;
  assign cache_tag__T_204_mask = 1'h0;
  assign cache_tag__T_204_en = reset;
  assign cache_tag__T_205_data = 24'h0;
  assign cache_tag__T_205_addr = 8'hc3;
  assign cache_tag__T_205_mask = 1'h0;
  assign cache_tag__T_205_en = reset;
  assign cache_tag__T_206_data = 24'h0;
  assign cache_tag__T_206_addr = 8'hc4;
  assign cache_tag__T_206_mask = 1'h0;
  assign cache_tag__T_206_en = reset;
  assign cache_tag__T_207_data = 24'h0;
  assign cache_tag__T_207_addr = 8'hc5;
  assign cache_tag__T_207_mask = 1'h0;
  assign cache_tag__T_207_en = reset;
  assign cache_tag__T_208_data = 24'h0;
  assign cache_tag__T_208_addr = 8'hc6;
  assign cache_tag__T_208_mask = 1'h0;
  assign cache_tag__T_208_en = reset;
  assign cache_tag__T_209_data = 24'h0;
  assign cache_tag__T_209_addr = 8'hc7;
  assign cache_tag__T_209_mask = 1'h0;
  assign cache_tag__T_209_en = reset;
  assign cache_tag__T_210_data = 24'h0;
  assign cache_tag__T_210_addr = 8'hc8;
  assign cache_tag__T_210_mask = 1'h0;
  assign cache_tag__T_210_en = reset;
  assign cache_tag__T_211_data = 24'h0;
  assign cache_tag__T_211_addr = 8'hc9;
  assign cache_tag__T_211_mask = 1'h0;
  assign cache_tag__T_211_en = reset;
  assign cache_tag__T_212_data = 24'h0;
  assign cache_tag__T_212_addr = 8'hca;
  assign cache_tag__T_212_mask = 1'h0;
  assign cache_tag__T_212_en = reset;
  assign cache_tag__T_213_data = 24'h0;
  assign cache_tag__T_213_addr = 8'hcb;
  assign cache_tag__T_213_mask = 1'h0;
  assign cache_tag__T_213_en = reset;
  assign cache_tag__T_214_data = 24'h0;
  assign cache_tag__T_214_addr = 8'hcc;
  assign cache_tag__T_214_mask = 1'h0;
  assign cache_tag__T_214_en = reset;
  assign cache_tag__T_215_data = 24'h0;
  assign cache_tag__T_215_addr = 8'hcd;
  assign cache_tag__T_215_mask = 1'h0;
  assign cache_tag__T_215_en = reset;
  assign cache_tag__T_216_data = 24'h0;
  assign cache_tag__T_216_addr = 8'hce;
  assign cache_tag__T_216_mask = 1'h0;
  assign cache_tag__T_216_en = reset;
  assign cache_tag__T_217_data = 24'h0;
  assign cache_tag__T_217_addr = 8'hcf;
  assign cache_tag__T_217_mask = 1'h0;
  assign cache_tag__T_217_en = reset;
  assign cache_tag__T_218_data = 24'h0;
  assign cache_tag__T_218_addr = 8'hd0;
  assign cache_tag__T_218_mask = 1'h0;
  assign cache_tag__T_218_en = reset;
  assign cache_tag__T_219_data = 24'h0;
  assign cache_tag__T_219_addr = 8'hd1;
  assign cache_tag__T_219_mask = 1'h0;
  assign cache_tag__T_219_en = reset;
  assign cache_tag__T_220_data = 24'h0;
  assign cache_tag__T_220_addr = 8'hd2;
  assign cache_tag__T_220_mask = 1'h0;
  assign cache_tag__T_220_en = reset;
  assign cache_tag__T_221_data = 24'h0;
  assign cache_tag__T_221_addr = 8'hd3;
  assign cache_tag__T_221_mask = 1'h0;
  assign cache_tag__T_221_en = reset;
  assign cache_tag__T_222_data = 24'h0;
  assign cache_tag__T_222_addr = 8'hd4;
  assign cache_tag__T_222_mask = 1'h0;
  assign cache_tag__T_222_en = reset;
  assign cache_tag__T_223_data = 24'h0;
  assign cache_tag__T_223_addr = 8'hd5;
  assign cache_tag__T_223_mask = 1'h0;
  assign cache_tag__T_223_en = reset;
  assign cache_tag__T_224_data = 24'h0;
  assign cache_tag__T_224_addr = 8'hd6;
  assign cache_tag__T_224_mask = 1'h0;
  assign cache_tag__T_224_en = reset;
  assign cache_tag__T_225_data = 24'h0;
  assign cache_tag__T_225_addr = 8'hd7;
  assign cache_tag__T_225_mask = 1'h0;
  assign cache_tag__T_225_en = reset;
  assign cache_tag__T_226_data = 24'h0;
  assign cache_tag__T_226_addr = 8'hd8;
  assign cache_tag__T_226_mask = 1'h0;
  assign cache_tag__T_226_en = reset;
  assign cache_tag__T_227_data = 24'h0;
  assign cache_tag__T_227_addr = 8'hd9;
  assign cache_tag__T_227_mask = 1'h0;
  assign cache_tag__T_227_en = reset;
  assign cache_tag__T_228_data = 24'h0;
  assign cache_tag__T_228_addr = 8'hda;
  assign cache_tag__T_228_mask = 1'h0;
  assign cache_tag__T_228_en = reset;
  assign cache_tag__T_229_data = 24'h0;
  assign cache_tag__T_229_addr = 8'hdb;
  assign cache_tag__T_229_mask = 1'h0;
  assign cache_tag__T_229_en = reset;
  assign cache_tag__T_230_data = 24'h0;
  assign cache_tag__T_230_addr = 8'hdc;
  assign cache_tag__T_230_mask = 1'h0;
  assign cache_tag__T_230_en = reset;
  assign cache_tag__T_231_data = 24'h0;
  assign cache_tag__T_231_addr = 8'hdd;
  assign cache_tag__T_231_mask = 1'h0;
  assign cache_tag__T_231_en = reset;
  assign cache_tag__T_232_data = 24'h0;
  assign cache_tag__T_232_addr = 8'hde;
  assign cache_tag__T_232_mask = 1'h0;
  assign cache_tag__T_232_en = reset;
  assign cache_tag__T_233_data = 24'h0;
  assign cache_tag__T_233_addr = 8'hdf;
  assign cache_tag__T_233_mask = 1'h0;
  assign cache_tag__T_233_en = reset;
  assign cache_tag__T_234_data = 24'h0;
  assign cache_tag__T_234_addr = 8'he0;
  assign cache_tag__T_234_mask = 1'h0;
  assign cache_tag__T_234_en = reset;
  assign cache_tag__T_235_data = 24'h0;
  assign cache_tag__T_235_addr = 8'he1;
  assign cache_tag__T_235_mask = 1'h0;
  assign cache_tag__T_235_en = reset;
  assign cache_tag__T_236_data = 24'h0;
  assign cache_tag__T_236_addr = 8'he2;
  assign cache_tag__T_236_mask = 1'h0;
  assign cache_tag__T_236_en = reset;
  assign cache_tag__T_237_data = 24'h0;
  assign cache_tag__T_237_addr = 8'he3;
  assign cache_tag__T_237_mask = 1'h0;
  assign cache_tag__T_237_en = reset;
  assign cache_tag__T_238_data = 24'h0;
  assign cache_tag__T_238_addr = 8'he4;
  assign cache_tag__T_238_mask = 1'h0;
  assign cache_tag__T_238_en = reset;
  assign cache_tag__T_239_data = 24'h0;
  assign cache_tag__T_239_addr = 8'he5;
  assign cache_tag__T_239_mask = 1'h0;
  assign cache_tag__T_239_en = reset;
  assign cache_tag__T_240_data = 24'h0;
  assign cache_tag__T_240_addr = 8'he6;
  assign cache_tag__T_240_mask = 1'h0;
  assign cache_tag__T_240_en = reset;
  assign cache_tag__T_241_data = 24'h0;
  assign cache_tag__T_241_addr = 8'he7;
  assign cache_tag__T_241_mask = 1'h0;
  assign cache_tag__T_241_en = reset;
  assign cache_tag__T_242_data = 24'h0;
  assign cache_tag__T_242_addr = 8'he8;
  assign cache_tag__T_242_mask = 1'h0;
  assign cache_tag__T_242_en = reset;
  assign cache_tag__T_243_data = 24'h0;
  assign cache_tag__T_243_addr = 8'he9;
  assign cache_tag__T_243_mask = 1'h0;
  assign cache_tag__T_243_en = reset;
  assign cache_tag__T_244_data = 24'h0;
  assign cache_tag__T_244_addr = 8'hea;
  assign cache_tag__T_244_mask = 1'h0;
  assign cache_tag__T_244_en = reset;
  assign cache_tag__T_245_data = 24'h0;
  assign cache_tag__T_245_addr = 8'heb;
  assign cache_tag__T_245_mask = 1'h0;
  assign cache_tag__T_245_en = reset;
  assign cache_tag__T_246_data = 24'h0;
  assign cache_tag__T_246_addr = 8'hec;
  assign cache_tag__T_246_mask = 1'h0;
  assign cache_tag__T_246_en = reset;
  assign cache_tag__T_247_data = 24'h0;
  assign cache_tag__T_247_addr = 8'hed;
  assign cache_tag__T_247_mask = 1'h0;
  assign cache_tag__T_247_en = reset;
  assign cache_tag__T_248_data = 24'h0;
  assign cache_tag__T_248_addr = 8'hee;
  assign cache_tag__T_248_mask = 1'h0;
  assign cache_tag__T_248_en = reset;
  assign cache_tag__T_249_data = 24'h0;
  assign cache_tag__T_249_addr = 8'hef;
  assign cache_tag__T_249_mask = 1'h0;
  assign cache_tag__T_249_en = reset;
  assign cache_tag__T_250_data = 24'h0;
  assign cache_tag__T_250_addr = 8'hf0;
  assign cache_tag__T_250_mask = 1'h0;
  assign cache_tag__T_250_en = reset;
  assign cache_tag__T_251_data = 24'h0;
  assign cache_tag__T_251_addr = 8'hf1;
  assign cache_tag__T_251_mask = 1'h0;
  assign cache_tag__T_251_en = reset;
  assign cache_tag__T_252_data = 24'h0;
  assign cache_tag__T_252_addr = 8'hf2;
  assign cache_tag__T_252_mask = 1'h0;
  assign cache_tag__T_252_en = reset;
  assign cache_tag__T_253_data = 24'h0;
  assign cache_tag__T_253_addr = 8'hf3;
  assign cache_tag__T_253_mask = 1'h0;
  assign cache_tag__T_253_en = reset;
  assign cache_tag__T_254_data = 24'h0;
  assign cache_tag__T_254_addr = 8'hf4;
  assign cache_tag__T_254_mask = 1'h0;
  assign cache_tag__T_254_en = reset;
  assign cache_tag__T_255_data = 24'h0;
  assign cache_tag__T_255_addr = 8'hf5;
  assign cache_tag__T_255_mask = 1'h0;
  assign cache_tag__T_255_en = reset;
  assign cache_tag__T_256_data = 24'h0;
  assign cache_tag__T_256_addr = 8'hf6;
  assign cache_tag__T_256_mask = 1'h0;
  assign cache_tag__T_256_en = reset;
  assign cache_tag__T_257_data = 24'h0;
  assign cache_tag__T_257_addr = 8'hf7;
  assign cache_tag__T_257_mask = 1'h0;
  assign cache_tag__T_257_en = reset;
  assign cache_tag__T_258_data = 24'h0;
  assign cache_tag__T_258_addr = 8'hf8;
  assign cache_tag__T_258_mask = 1'h0;
  assign cache_tag__T_258_en = reset;
  assign cache_tag__T_259_data = 24'h0;
  assign cache_tag__T_259_addr = 8'hf9;
  assign cache_tag__T_259_mask = 1'h0;
  assign cache_tag__T_259_en = reset;
  assign cache_tag__T_260_data = 24'h0;
  assign cache_tag__T_260_addr = 8'hfa;
  assign cache_tag__T_260_mask = 1'h0;
  assign cache_tag__T_260_en = reset;
  assign cache_tag__T_261_data = 24'h0;
  assign cache_tag__T_261_addr = 8'hfb;
  assign cache_tag__T_261_mask = 1'h0;
  assign cache_tag__T_261_en = reset;
  assign cache_tag__T_262_data = 24'h0;
  assign cache_tag__T_262_addr = 8'hfc;
  assign cache_tag__T_262_mask = 1'h0;
  assign cache_tag__T_262_en = reset;
  assign cache_tag__T_263_data = 24'h0;
  assign cache_tag__T_263_addr = 8'hfd;
  assign cache_tag__T_263_mask = 1'h0;
  assign cache_tag__T_263_en = reset;
  assign cache_tag__T_264_data = 24'h0;
  assign cache_tag__T_264_addr = 8'hfe;
  assign cache_tag__T_264_mask = 1'h0;
  assign cache_tag__T_264_en = reset;
  assign cache_tag__T_265_data = 24'h0;
  assign cache_tag__T_265_addr = 8'hff;
  assign cache_tag__T_265_mask = 1'h0;
  assign cache_tag__T_265_en = reset;
  assign cache_tag_s1_entry_w_data = s1_in_addr[31:8];
  assign cache_tag_s1_entry_w_addr = s1_in_addr[7:0];
  assign cache_tag_s1_entry_w_mask = s1_resp & _T_285;
  assign cache_tag_s1_entry_w_en = s1_resp & _T_285;
  assign cache_data_s1_entry_r_addr = s1_in_addr[7:0];
  assign cache_data_s1_entry_r_data = cache_data[cache_data_s1_entry_r_addr]; // @[icache.scala 91:18]
  assign cache_data__T_8_data = 32'h0;
  assign cache_data__T_8_addr = _T_6[7:0];
  assign cache_data__T_8_mask = 1'h0;
  assign cache_data__T_8_en = _T_1 & _T_5;
  assign cache_data__T_10_data = 32'h0;
  assign cache_data__T_10_addr = 8'h0;
  assign cache_data__T_10_mask = 1'h0;
  assign cache_data__T_10_en = reset;
  assign cache_data__T_11_data = 32'h0;
  assign cache_data__T_11_addr = 8'h1;
  assign cache_data__T_11_mask = 1'h0;
  assign cache_data__T_11_en = reset;
  assign cache_data__T_12_data = 32'h0;
  assign cache_data__T_12_addr = 8'h2;
  assign cache_data__T_12_mask = 1'h0;
  assign cache_data__T_12_en = reset;
  assign cache_data__T_13_data = 32'h0;
  assign cache_data__T_13_addr = 8'h3;
  assign cache_data__T_13_mask = 1'h0;
  assign cache_data__T_13_en = reset;
  assign cache_data__T_14_data = 32'h0;
  assign cache_data__T_14_addr = 8'h4;
  assign cache_data__T_14_mask = 1'h0;
  assign cache_data__T_14_en = reset;
  assign cache_data__T_15_data = 32'h0;
  assign cache_data__T_15_addr = 8'h5;
  assign cache_data__T_15_mask = 1'h0;
  assign cache_data__T_15_en = reset;
  assign cache_data__T_16_data = 32'h0;
  assign cache_data__T_16_addr = 8'h6;
  assign cache_data__T_16_mask = 1'h0;
  assign cache_data__T_16_en = reset;
  assign cache_data__T_17_data = 32'h0;
  assign cache_data__T_17_addr = 8'h7;
  assign cache_data__T_17_mask = 1'h0;
  assign cache_data__T_17_en = reset;
  assign cache_data__T_18_data = 32'h0;
  assign cache_data__T_18_addr = 8'h8;
  assign cache_data__T_18_mask = 1'h0;
  assign cache_data__T_18_en = reset;
  assign cache_data__T_19_data = 32'h0;
  assign cache_data__T_19_addr = 8'h9;
  assign cache_data__T_19_mask = 1'h0;
  assign cache_data__T_19_en = reset;
  assign cache_data__T_20_data = 32'h0;
  assign cache_data__T_20_addr = 8'ha;
  assign cache_data__T_20_mask = 1'h0;
  assign cache_data__T_20_en = reset;
  assign cache_data__T_21_data = 32'h0;
  assign cache_data__T_21_addr = 8'hb;
  assign cache_data__T_21_mask = 1'h0;
  assign cache_data__T_21_en = reset;
  assign cache_data__T_22_data = 32'h0;
  assign cache_data__T_22_addr = 8'hc;
  assign cache_data__T_22_mask = 1'h0;
  assign cache_data__T_22_en = reset;
  assign cache_data__T_23_data = 32'h0;
  assign cache_data__T_23_addr = 8'hd;
  assign cache_data__T_23_mask = 1'h0;
  assign cache_data__T_23_en = reset;
  assign cache_data__T_24_data = 32'h0;
  assign cache_data__T_24_addr = 8'he;
  assign cache_data__T_24_mask = 1'h0;
  assign cache_data__T_24_en = reset;
  assign cache_data__T_25_data = 32'h0;
  assign cache_data__T_25_addr = 8'hf;
  assign cache_data__T_25_mask = 1'h0;
  assign cache_data__T_25_en = reset;
  assign cache_data__T_26_data = 32'h0;
  assign cache_data__T_26_addr = 8'h10;
  assign cache_data__T_26_mask = 1'h0;
  assign cache_data__T_26_en = reset;
  assign cache_data__T_27_data = 32'h0;
  assign cache_data__T_27_addr = 8'h11;
  assign cache_data__T_27_mask = 1'h0;
  assign cache_data__T_27_en = reset;
  assign cache_data__T_28_data = 32'h0;
  assign cache_data__T_28_addr = 8'h12;
  assign cache_data__T_28_mask = 1'h0;
  assign cache_data__T_28_en = reset;
  assign cache_data__T_29_data = 32'h0;
  assign cache_data__T_29_addr = 8'h13;
  assign cache_data__T_29_mask = 1'h0;
  assign cache_data__T_29_en = reset;
  assign cache_data__T_30_data = 32'h0;
  assign cache_data__T_30_addr = 8'h14;
  assign cache_data__T_30_mask = 1'h0;
  assign cache_data__T_30_en = reset;
  assign cache_data__T_31_data = 32'h0;
  assign cache_data__T_31_addr = 8'h15;
  assign cache_data__T_31_mask = 1'h0;
  assign cache_data__T_31_en = reset;
  assign cache_data__T_32_data = 32'h0;
  assign cache_data__T_32_addr = 8'h16;
  assign cache_data__T_32_mask = 1'h0;
  assign cache_data__T_32_en = reset;
  assign cache_data__T_33_data = 32'h0;
  assign cache_data__T_33_addr = 8'h17;
  assign cache_data__T_33_mask = 1'h0;
  assign cache_data__T_33_en = reset;
  assign cache_data__T_34_data = 32'h0;
  assign cache_data__T_34_addr = 8'h18;
  assign cache_data__T_34_mask = 1'h0;
  assign cache_data__T_34_en = reset;
  assign cache_data__T_35_data = 32'h0;
  assign cache_data__T_35_addr = 8'h19;
  assign cache_data__T_35_mask = 1'h0;
  assign cache_data__T_35_en = reset;
  assign cache_data__T_36_data = 32'h0;
  assign cache_data__T_36_addr = 8'h1a;
  assign cache_data__T_36_mask = 1'h0;
  assign cache_data__T_36_en = reset;
  assign cache_data__T_37_data = 32'h0;
  assign cache_data__T_37_addr = 8'h1b;
  assign cache_data__T_37_mask = 1'h0;
  assign cache_data__T_37_en = reset;
  assign cache_data__T_38_data = 32'h0;
  assign cache_data__T_38_addr = 8'h1c;
  assign cache_data__T_38_mask = 1'h0;
  assign cache_data__T_38_en = reset;
  assign cache_data__T_39_data = 32'h0;
  assign cache_data__T_39_addr = 8'h1d;
  assign cache_data__T_39_mask = 1'h0;
  assign cache_data__T_39_en = reset;
  assign cache_data__T_40_data = 32'h0;
  assign cache_data__T_40_addr = 8'h1e;
  assign cache_data__T_40_mask = 1'h0;
  assign cache_data__T_40_en = reset;
  assign cache_data__T_41_data = 32'h0;
  assign cache_data__T_41_addr = 8'h1f;
  assign cache_data__T_41_mask = 1'h0;
  assign cache_data__T_41_en = reset;
  assign cache_data__T_42_data = 32'h0;
  assign cache_data__T_42_addr = 8'h20;
  assign cache_data__T_42_mask = 1'h0;
  assign cache_data__T_42_en = reset;
  assign cache_data__T_43_data = 32'h0;
  assign cache_data__T_43_addr = 8'h21;
  assign cache_data__T_43_mask = 1'h0;
  assign cache_data__T_43_en = reset;
  assign cache_data__T_44_data = 32'h0;
  assign cache_data__T_44_addr = 8'h22;
  assign cache_data__T_44_mask = 1'h0;
  assign cache_data__T_44_en = reset;
  assign cache_data__T_45_data = 32'h0;
  assign cache_data__T_45_addr = 8'h23;
  assign cache_data__T_45_mask = 1'h0;
  assign cache_data__T_45_en = reset;
  assign cache_data__T_46_data = 32'h0;
  assign cache_data__T_46_addr = 8'h24;
  assign cache_data__T_46_mask = 1'h0;
  assign cache_data__T_46_en = reset;
  assign cache_data__T_47_data = 32'h0;
  assign cache_data__T_47_addr = 8'h25;
  assign cache_data__T_47_mask = 1'h0;
  assign cache_data__T_47_en = reset;
  assign cache_data__T_48_data = 32'h0;
  assign cache_data__T_48_addr = 8'h26;
  assign cache_data__T_48_mask = 1'h0;
  assign cache_data__T_48_en = reset;
  assign cache_data__T_49_data = 32'h0;
  assign cache_data__T_49_addr = 8'h27;
  assign cache_data__T_49_mask = 1'h0;
  assign cache_data__T_49_en = reset;
  assign cache_data__T_50_data = 32'h0;
  assign cache_data__T_50_addr = 8'h28;
  assign cache_data__T_50_mask = 1'h0;
  assign cache_data__T_50_en = reset;
  assign cache_data__T_51_data = 32'h0;
  assign cache_data__T_51_addr = 8'h29;
  assign cache_data__T_51_mask = 1'h0;
  assign cache_data__T_51_en = reset;
  assign cache_data__T_52_data = 32'h0;
  assign cache_data__T_52_addr = 8'h2a;
  assign cache_data__T_52_mask = 1'h0;
  assign cache_data__T_52_en = reset;
  assign cache_data__T_53_data = 32'h0;
  assign cache_data__T_53_addr = 8'h2b;
  assign cache_data__T_53_mask = 1'h0;
  assign cache_data__T_53_en = reset;
  assign cache_data__T_54_data = 32'h0;
  assign cache_data__T_54_addr = 8'h2c;
  assign cache_data__T_54_mask = 1'h0;
  assign cache_data__T_54_en = reset;
  assign cache_data__T_55_data = 32'h0;
  assign cache_data__T_55_addr = 8'h2d;
  assign cache_data__T_55_mask = 1'h0;
  assign cache_data__T_55_en = reset;
  assign cache_data__T_56_data = 32'h0;
  assign cache_data__T_56_addr = 8'h2e;
  assign cache_data__T_56_mask = 1'h0;
  assign cache_data__T_56_en = reset;
  assign cache_data__T_57_data = 32'h0;
  assign cache_data__T_57_addr = 8'h2f;
  assign cache_data__T_57_mask = 1'h0;
  assign cache_data__T_57_en = reset;
  assign cache_data__T_58_data = 32'h0;
  assign cache_data__T_58_addr = 8'h30;
  assign cache_data__T_58_mask = 1'h0;
  assign cache_data__T_58_en = reset;
  assign cache_data__T_59_data = 32'h0;
  assign cache_data__T_59_addr = 8'h31;
  assign cache_data__T_59_mask = 1'h0;
  assign cache_data__T_59_en = reset;
  assign cache_data__T_60_data = 32'h0;
  assign cache_data__T_60_addr = 8'h32;
  assign cache_data__T_60_mask = 1'h0;
  assign cache_data__T_60_en = reset;
  assign cache_data__T_61_data = 32'h0;
  assign cache_data__T_61_addr = 8'h33;
  assign cache_data__T_61_mask = 1'h0;
  assign cache_data__T_61_en = reset;
  assign cache_data__T_62_data = 32'h0;
  assign cache_data__T_62_addr = 8'h34;
  assign cache_data__T_62_mask = 1'h0;
  assign cache_data__T_62_en = reset;
  assign cache_data__T_63_data = 32'h0;
  assign cache_data__T_63_addr = 8'h35;
  assign cache_data__T_63_mask = 1'h0;
  assign cache_data__T_63_en = reset;
  assign cache_data__T_64_data = 32'h0;
  assign cache_data__T_64_addr = 8'h36;
  assign cache_data__T_64_mask = 1'h0;
  assign cache_data__T_64_en = reset;
  assign cache_data__T_65_data = 32'h0;
  assign cache_data__T_65_addr = 8'h37;
  assign cache_data__T_65_mask = 1'h0;
  assign cache_data__T_65_en = reset;
  assign cache_data__T_66_data = 32'h0;
  assign cache_data__T_66_addr = 8'h38;
  assign cache_data__T_66_mask = 1'h0;
  assign cache_data__T_66_en = reset;
  assign cache_data__T_67_data = 32'h0;
  assign cache_data__T_67_addr = 8'h39;
  assign cache_data__T_67_mask = 1'h0;
  assign cache_data__T_67_en = reset;
  assign cache_data__T_68_data = 32'h0;
  assign cache_data__T_68_addr = 8'h3a;
  assign cache_data__T_68_mask = 1'h0;
  assign cache_data__T_68_en = reset;
  assign cache_data__T_69_data = 32'h0;
  assign cache_data__T_69_addr = 8'h3b;
  assign cache_data__T_69_mask = 1'h0;
  assign cache_data__T_69_en = reset;
  assign cache_data__T_70_data = 32'h0;
  assign cache_data__T_70_addr = 8'h3c;
  assign cache_data__T_70_mask = 1'h0;
  assign cache_data__T_70_en = reset;
  assign cache_data__T_71_data = 32'h0;
  assign cache_data__T_71_addr = 8'h3d;
  assign cache_data__T_71_mask = 1'h0;
  assign cache_data__T_71_en = reset;
  assign cache_data__T_72_data = 32'h0;
  assign cache_data__T_72_addr = 8'h3e;
  assign cache_data__T_72_mask = 1'h0;
  assign cache_data__T_72_en = reset;
  assign cache_data__T_73_data = 32'h0;
  assign cache_data__T_73_addr = 8'h3f;
  assign cache_data__T_73_mask = 1'h0;
  assign cache_data__T_73_en = reset;
  assign cache_data__T_74_data = 32'h0;
  assign cache_data__T_74_addr = 8'h40;
  assign cache_data__T_74_mask = 1'h0;
  assign cache_data__T_74_en = reset;
  assign cache_data__T_75_data = 32'h0;
  assign cache_data__T_75_addr = 8'h41;
  assign cache_data__T_75_mask = 1'h0;
  assign cache_data__T_75_en = reset;
  assign cache_data__T_76_data = 32'h0;
  assign cache_data__T_76_addr = 8'h42;
  assign cache_data__T_76_mask = 1'h0;
  assign cache_data__T_76_en = reset;
  assign cache_data__T_77_data = 32'h0;
  assign cache_data__T_77_addr = 8'h43;
  assign cache_data__T_77_mask = 1'h0;
  assign cache_data__T_77_en = reset;
  assign cache_data__T_78_data = 32'h0;
  assign cache_data__T_78_addr = 8'h44;
  assign cache_data__T_78_mask = 1'h0;
  assign cache_data__T_78_en = reset;
  assign cache_data__T_79_data = 32'h0;
  assign cache_data__T_79_addr = 8'h45;
  assign cache_data__T_79_mask = 1'h0;
  assign cache_data__T_79_en = reset;
  assign cache_data__T_80_data = 32'h0;
  assign cache_data__T_80_addr = 8'h46;
  assign cache_data__T_80_mask = 1'h0;
  assign cache_data__T_80_en = reset;
  assign cache_data__T_81_data = 32'h0;
  assign cache_data__T_81_addr = 8'h47;
  assign cache_data__T_81_mask = 1'h0;
  assign cache_data__T_81_en = reset;
  assign cache_data__T_82_data = 32'h0;
  assign cache_data__T_82_addr = 8'h48;
  assign cache_data__T_82_mask = 1'h0;
  assign cache_data__T_82_en = reset;
  assign cache_data__T_83_data = 32'h0;
  assign cache_data__T_83_addr = 8'h49;
  assign cache_data__T_83_mask = 1'h0;
  assign cache_data__T_83_en = reset;
  assign cache_data__T_84_data = 32'h0;
  assign cache_data__T_84_addr = 8'h4a;
  assign cache_data__T_84_mask = 1'h0;
  assign cache_data__T_84_en = reset;
  assign cache_data__T_85_data = 32'h0;
  assign cache_data__T_85_addr = 8'h4b;
  assign cache_data__T_85_mask = 1'h0;
  assign cache_data__T_85_en = reset;
  assign cache_data__T_86_data = 32'h0;
  assign cache_data__T_86_addr = 8'h4c;
  assign cache_data__T_86_mask = 1'h0;
  assign cache_data__T_86_en = reset;
  assign cache_data__T_87_data = 32'h0;
  assign cache_data__T_87_addr = 8'h4d;
  assign cache_data__T_87_mask = 1'h0;
  assign cache_data__T_87_en = reset;
  assign cache_data__T_88_data = 32'h0;
  assign cache_data__T_88_addr = 8'h4e;
  assign cache_data__T_88_mask = 1'h0;
  assign cache_data__T_88_en = reset;
  assign cache_data__T_89_data = 32'h0;
  assign cache_data__T_89_addr = 8'h4f;
  assign cache_data__T_89_mask = 1'h0;
  assign cache_data__T_89_en = reset;
  assign cache_data__T_90_data = 32'h0;
  assign cache_data__T_90_addr = 8'h50;
  assign cache_data__T_90_mask = 1'h0;
  assign cache_data__T_90_en = reset;
  assign cache_data__T_91_data = 32'h0;
  assign cache_data__T_91_addr = 8'h51;
  assign cache_data__T_91_mask = 1'h0;
  assign cache_data__T_91_en = reset;
  assign cache_data__T_92_data = 32'h0;
  assign cache_data__T_92_addr = 8'h52;
  assign cache_data__T_92_mask = 1'h0;
  assign cache_data__T_92_en = reset;
  assign cache_data__T_93_data = 32'h0;
  assign cache_data__T_93_addr = 8'h53;
  assign cache_data__T_93_mask = 1'h0;
  assign cache_data__T_93_en = reset;
  assign cache_data__T_94_data = 32'h0;
  assign cache_data__T_94_addr = 8'h54;
  assign cache_data__T_94_mask = 1'h0;
  assign cache_data__T_94_en = reset;
  assign cache_data__T_95_data = 32'h0;
  assign cache_data__T_95_addr = 8'h55;
  assign cache_data__T_95_mask = 1'h0;
  assign cache_data__T_95_en = reset;
  assign cache_data__T_96_data = 32'h0;
  assign cache_data__T_96_addr = 8'h56;
  assign cache_data__T_96_mask = 1'h0;
  assign cache_data__T_96_en = reset;
  assign cache_data__T_97_data = 32'h0;
  assign cache_data__T_97_addr = 8'h57;
  assign cache_data__T_97_mask = 1'h0;
  assign cache_data__T_97_en = reset;
  assign cache_data__T_98_data = 32'h0;
  assign cache_data__T_98_addr = 8'h58;
  assign cache_data__T_98_mask = 1'h0;
  assign cache_data__T_98_en = reset;
  assign cache_data__T_99_data = 32'h0;
  assign cache_data__T_99_addr = 8'h59;
  assign cache_data__T_99_mask = 1'h0;
  assign cache_data__T_99_en = reset;
  assign cache_data__T_100_data = 32'h0;
  assign cache_data__T_100_addr = 8'h5a;
  assign cache_data__T_100_mask = 1'h0;
  assign cache_data__T_100_en = reset;
  assign cache_data__T_101_data = 32'h0;
  assign cache_data__T_101_addr = 8'h5b;
  assign cache_data__T_101_mask = 1'h0;
  assign cache_data__T_101_en = reset;
  assign cache_data__T_102_data = 32'h0;
  assign cache_data__T_102_addr = 8'h5c;
  assign cache_data__T_102_mask = 1'h0;
  assign cache_data__T_102_en = reset;
  assign cache_data__T_103_data = 32'h0;
  assign cache_data__T_103_addr = 8'h5d;
  assign cache_data__T_103_mask = 1'h0;
  assign cache_data__T_103_en = reset;
  assign cache_data__T_104_data = 32'h0;
  assign cache_data__T_104_addr = 8'h5e;
  assign cache_data__T_104_mask = 1'h0;
  assign cache_data__T_104_en = reset;
  assign cache_data__T_105_data = 32'h0;
  assign cache_data__T_105_addr = 8'h5f;
  assign cache_data__T_105_mask = 1'h0;
  assign cache_data__T_105_en = reset;
  assign cache_data__T_106_data = 32'h0;
  assign cache_data__T_106_addr = 8'h60;
  assign cache_data__T_106_mask = 1'h0;
  assign cache_data__T_106_en = reset;
  assign cache_data__T_107_data = 32'h0;
  assign cache_data__T_107_addr = 8'h61;
  assign cache_data__T_107_mask = 1'h0;
  assign cache_data__T_107_en = reset;
  assign cache_data__T_108_data = 32'h0;
  assign cache_data__T_108_addr = 8'h62;
  assign cache_data__T_108_mask = 1'h0;
  assign cache_data__T_108_en = reset;
  assign cache_data__T_109_data = 32'h0;
  assign cache_data__T_109_addr = 8'h63;
  assign cache_data__T_109_mask = 1'h0;
  assign cache_data__T_109_en = reset;
  assign cache_data__T_110_data = 32'h0;
  assign cache_data__T_110_addr = 8'h64;
  assign cache_data__T_110_mask = 1'h0;
  assign cache_data__T_110_en = reset;
  assign cache_data__T_111_data = 32'h0;
  assign cache_data__T_111_addr = 8'h65;
  assign cache_data__T_111_mask = 1'h0;
  assign cache_data__T_111_en = reset;
  assign cache_data__T_112_data = 32'h0;
  assign cache_data__T_112_addr = 8'h66;
  assign cache_data__T_112_mask = 1'h0;
  assign cache_data__T_112_en = reset;
  assign cache_data__T_113_data = 32'h0;
  assign cache_data__T_113_addr = 8'h67;
  assign cache_data__T_113_mask = 1'h0;
  assign cache_data__T_113_en = reset;
  assign cache_data__T_114_data = 32'h0;
  assign cache_data__T_114_addr = 8'h68;
  assign cache_data__T_114_mask = 1'h0;
  assign cache_data__T_114_en = reset;
  assign cache_data__T_115_data = 32'h0;
  assign cache_data__T_115_addr = 8'h69;
  assign cache_data__T_115_mask = 1'h0;
  assign cache_data__T_115_en = reset;
  assign cache_data__T_116_data = 32'h0;
  assign cache_data__T_116_addr = 8'h6a;
  assign cache_data__T_116_mask = 1'h0;
  assign cache_data__T_116_en = reset;
  assign cache_data__T_117_data = 32'h0;
  assign cache_data__T_117_addr = 8'h6b;
  assign cache_data__T_117_mask = 1'h0;
  assign cache_data__T_117_en = reset;
  assign cache_data__T_118_data = 32'h0;
  assign cache_data__T_118_addr = 8'h6c;
  assign cache_data__T_118_mask = 1'h0;
  assign cache_data__T_118_en = reset;
  assign cache_data__T_119_data = 32'h0;
  assign cache_data__T_119_addr = 8'h6d;
  assign cache_data__T_119_mask = 1'h0;
  assign cache_data__T_119_en = reset;
  assign cache_data__T_120_data = 32'h0;
  assign cache_data__T_120_addr = 8'h6e;
  assign cache_data__T_120_mask = 1'h0;
  assign cache_data__T_120_en = reset;
  assign cache_data__T_121_data = 32'h0;
  assign cache_data__T_121_addr = 8'h6f;
  assign cache_data__T_121_mask = 1'h0;
  assign cache_data__T_121_en = reset;
  assign cache_data__T_122_data = 32'h0;
  assign cache_data__T_122_addr = 8'h70;
  assign cache_data__T_122_mask = 1'h0;
  assign cache_data__T_122_en = reset;
  assign cache_data__T_123_data = 32'h0;
  assign cache_data__T_123_addr = 8'h71;
  assign cache_data__T_123_mask = 1'h0;
  assign cache_data__T_123_en = reset;
  assign cache_data__T_124_data = 32'h0;
  assign cache_data__T_124_addr = 8'h72;
  assign cache_data__T_124_mask = 1'h0;
  assign cache_data__T_124_en = reset;
  assign cache_data__T_125_data = 32'h0;
  assign cache_data__T_125_addr = 8'h73;
  assign cache_data__T_125_mask = 1'h0;
  assign cache_data__T_125_en = reset;
  assign cache_data__T_126_data = 32'h0;
  assign cache_data__T_126_addr = 8'h74;
  assign cache_data__T_126_mask = 1'h0;
  assign cache_data__T_126_en = reset;
  assign cache_data__T_127_data = 32'h0;
  assign cache_data__T_127_addr = 8'h75;
  assign cache_data__T_127_mask = 1'h0;
  assign cache_data__T_127_en = reset;
  assign cache_data__T_128_data = 32'h0;
  assign cache_data__T_128_addr = 8'h76;
  assign cache_data__T_128_mask = 1'h0;
  assign cache_data__T_128_en = reset;
  assign cache_data__T_129_data = 32'h0;
  assign cache_data__T_129_addr = 8'h77;
  assign cache_data__T_129_mask = 1'h0;
  assign cache_data__T_129_en = reset;
  assign cache_data__T_130_data = 32'h0;
  assign cache_data__T_130_addr = 8'h78;
  assign cache_data__T_130_mask = 1'h0;
  assign cache_data__T_130_en = reset;
  assign cache_data__T_131_data = 32'h0;
  assign cache_data__T_131_addr = 8'h79;
  assign cache_data__T_131_mask = 1'h0;
  assign cache_data__T_131_en = reset;
  assign cache_data__T_132_data = 32'h0;
  assign cache_data__T_132_addr = 8'h7a;
  assign cache_data__T_132_mask = 1'h0;
  assign cache_data__T_132_en = reset;
  assign cache_data__T_133_data = 32'h0;
  assign cache_data__T_133_addr = 8'h7b;
  assign cache_data__T_133_mask = 1'h0;
  assign cache_data__T_133_en = reset;
  assign cache_data__T_134_data = 32'h0;
  assign cache_data__T_134_addr = 8'h7c;
  assign cache_data__T_134_mask = 1'h0;
  assign cache_data__T_134_en = reset;
  assign cache_data__T_135_data = 32'h0;
  assign cache_data__T_135_addr = 8'h7d;
  assign cache_data__T_135_mask = 1'h0;
  assign cache_data__T_135_en = reset;
  assign cache_data__T_136_data = 32'h0;
  assign cache_data__T_136_addr = 8'h7e;
  assign cache_data__T_136_mask = 1'h0;
  assign cache_data__T_136_en = reset;
  assign cache_data__T_137_data = 32'h0;
  assign cache_data__T_137_addr = 8'h7f;
  assign cache_data__T_137_mask = 1'h0;
  assign cache_data__T_137_en = reset;
  assign cache_data__T_138_data = 32'h0;
  assign cache_data__T_138_addr = 8'h80;
  assign cache_data__T_138_mask = 1'h0;
  assign cache_data__T_138_en = reset;
  assign cache_data__T_139_data = 32'h0;
  assign cache_data__T_139_addr = 8'h81;
  assign cache_data__T_139_mask = 1'h0;
  assign cache_data__T_139_en = reset;
  assign cache_data__T_140_data = 32'h0;
  assign cache_data__T_140_addr = 8'h82;
  assign cache_data__T_140_mask = 1'h0;
  assign cache_data__T_140_en = reset;
  assign cache_data__T_141_data = 32'h0;
  assign cache_data__T_141_addr = 8'h83;
  assign cache_data__T_141_mask = 1'h0;
  assign cache_data__T_141_en = reset;
  assign cache_data__T_142_data = 32'h0;
  assign cache_data__T_142_addr = 8'h84;
  assign cache_data__T_142_mask = 1'h0;
  assign cache_data__T_142_en = reset;
  assign cache_data__T_143_data = 32'h0;
  assign cache_data__T_143_addr = 8'h85;
  assign cache_data__T_143_mask = 1'h0;
  assign cache_data__T_143_en = reset;
  assign cache_data__T_144_data = 32'h0;
  assign cache_data__T_144_addr = 8'h86;
  assign cache_data__T_144_mask = 1'h0;
  assign cache_data__T_144_en = reset;
  assign cache_data__T_145_data = 32'h0;
  assign cache_data__T_145_addr = 8'h87;
  assign cache_data__T_145_mask = 1'h0;
  assign cache_data__T_145_en = reset;
  assign cache_data__T_146_data = 32'h0;
  assign cache_data__T_146_addr = 8'h88;
  assign cache_data__T_146_mask = 1'h0;
  assign cache_data__T_146_en = reset;
  assign cache_data__T_147_data = 32'h0;
  assign cache_data__T_147_addr = 8'h89;
  assign cache_data__T_147_mask = 1'h0;
  assign cache_data__T_147_en = reset;
  assign cache_data__T_148_data = 32'h0;
  assign cache_data__T_148_addr = 8'h8a;
  assign cache_data__T_148_mask = 1'h0;
  assign cache_data__T_148_en = reset;
  assign cache_data__T_149_data = 32'h0;
  assign cache_data__T_149_addr = 8'h8b;
  assign cache_data__T_149_mask = 1'h0;
  assign cache_data__T_149_en = reset;
  assign cache_data__T_150_data = 32'h0;
  assign cache_data__T_150_addr = 8'h8c;
  assign cache_data__T_150_mask = 1'h0;
  assign cache_data__T_150_en = reset;
  assign cache_data__T_151_data = 32'h0;
  assign cache_data__T_151_addr = 8'h8d;
  assign cache_data__T_151_mask = 1'h0;
  assign cache_data__T_151_en = reset;
  assign cache_data__T_152_data = 32'h0;
  assign cache_data__T_152_addr = 8'h8e;
  assign cache_data__T_152_mask = 1'h0;
  assign cache_data__T_152_en = reset;
  assign cache_data__T_153_data = 32'h0;
  assign cache_data__T_153_addr = 8'h8f;
  assign cache_data__T_153_mask = 1'h0;
  assign cache_data__T_153_en = reset;
  assign cache_data__T_154_data = 32'h0;
  assign cache_data__T_154_addr = 8'h90;
  assign cache_data__T_154_mask = 1'h0;
  assign cache_data__T_154_en = reset;
  assign cache_data__T_155_data = 32'h0;
  assign cache_data__T_155_addr = 8'h91;
  assign cache_data__T_155_mask = 1'h0;
  assign cache_data__T_155_en = reset;
  assign cache_data__T_156_data = 32'h0;
  assign cache_data__T_156_addr = 8'h92;
  assign cache_data__T_156_mask = 1'h0;
  assign cache_data__T_156_en = reset;
  assign cache_data__T_157_data = 32'h0;
  assign cache_data__T_157_addr = 8'h93;
  assign cache_data__T_157_mask = 1'h0;
  assign cache_data__T_157_en = reset;
  assign cache_data__T_158_data = 32'h0;
  assign cache_data__T_158_addr = 8'h94;
  assign cache_data__T_158_mask = 1'h0;
  assign cache_data__T_158_en = reset;
  assign cache_data__T_159_data = 32'h0;
  assign cache_data__T_159_addr = 8'h95;
  assign cache_data__T_159_mask = 1'h0;
  assign cache_data__T_159_en = reset;
  assign cache_data__T_160_data = 32'h0;
  assign cache_data__T_160_addr = 8'h96;
  assign cache_data__T_160_mask = 1'h0;
  assign cache_data__T_160_en = reset;
  assign cache_data__T_161_data = 32'h0;
  assign cache_data__T_161_addr = 8'h97;
  assign cache_data__T_161_mask = 1'h0;
  assign cache_data__T_161_en = reset;
  assign cache_data__T_162_data = 32'h0;
  assign cache_data__T_162_addr = 8'h98;
  assign cache_data__T_162_mask = 1'h0;
  assign cache_data__T_162_en = reset;
  assign cache_data__T_163_data = 32'h0;
  assign cache_data__T_163_addr = 8'h99;
  assign cache_data__T_163_mask = 1'h0;
  assign cache_data__T_163_en = reset;
  assign cache_data__T_164_data = 32'h0;
  assign cache_data__T_164_addr = 8'h9a;
  assign cache_data__T_164_mask = 1'h0;
  assign cache_data__T_164_en = reset;
  assign cache_data__T_165_data = 32'h0;
  assign cache_data__T_165_addr = 8'h9b;
  assign cache_data__T_165_mask = 1'h0;
  assign cache_data__T_165_en = reset;
  assign cache_data__T_166_data = 32'h0;
  assign cache_data__T_166_addr = 8'h9c;
  assign cache_data__T_166_mask = 1'h0;
  assign cache_data__T_166_en = reset;
  assign cache_data__T_167_data = 32'h0;
  assign cache_data__T_167_addr = 8'h9d;
  assign cache_data__T_167_mask = 1'h0;
  assign cache_data__T_167_en = reset;
  assign cache_data__T_168_data = 32'h0;
  assign cache_data__T_168_addr = 8'h9e;
  assign cache_data__T_168_mask = 1'h0;
  assign cache_data__T_168_en = reset;
  assign cache_data__T_169_data = 32'h0;
  assign cache_data__T_169_addr = 8'h9f;
  assign cache_data__T_169_mask = 1'h0;
  assign cache_data__T_169_en = reset;
  assign cache_data__T_170_data = 32'h0;
  assign cache_data__T_170_addr = 8'ha0;
  assign cache_data__T_170_mask = 1'h0;
  assign cache_data__T_170_en = reset;
  assign cache_data__T_171_data = 32'h0;
  assign cache_data__T_171_addr = 8'ha1;
  assign cache_data__T_171_mask = 1'h0;
  assign cache_data__T_171_en = reset;
  assign cache_data__T_172_data = 32'h0;
  assign cache_data__T_172_addr = 8'ha2;
  assign cache_data__T_172_mask = 1'h0;
  assign cache_data__T_172_en = reset;
  assign cache_data__T_173_data = 32'h0;
  assign cache_data__T_173_addr = 8'ha3;
  assign cache_data__T_173_mask = 1'h0;
  assign cache_data__T_173_en = reset;
  assign cache_data__T_174_data = 32'h0;
  assign cache_data__T_174_addr = 8'ha4;
  assign cache_data__T_174_mask = 1'h0;
  assign cache_data__T_174_en = reset;
  assign cache_data__T_175_data = 32'h0;
  assign cache_data__T_175_addr = 8'ha5;
  assign cache_data__T_175_mask = 1'h0;
  assign cache_data__T_175_en = reset;
  assign cache_data__T_176_data = 32'h0;
  assign cache_data__T_176_addr = 8'ha6;
  assign cache_data__T_176_mask = 1'h0;
  assign cache_data__T_176_en = reset;
  assign cache_data__T_177_data = 32'h0;
  assign cache_data__T_177_addr = 8'ha7;
  assign cache_data__T_177_mask = 1'h0;
  assign cache_data__T_177_en = reset;
  assign cache_data__T_178_data = 32'h0;
  assign cache_data__T_178_addr = 8'ha8;
  assign cache_data__T_178_mask = 1'h0;
  assign cache_data__T_178_en = reset;
  assign cache_data__T_179_data = 32'h0;
  assign cache_data__T_179_addr = 8'ha9;
  assign cache_data__T_179_mask = 1'h0;
  assign cache_data__T_179_en = reset;
  assign cache_data__T_180_data = 32'h0;
  assign cache_data__T_180_addr = 8'haa;
  assign cache_data__T_180_mask = 1'h0;
  assign cache_data__T_180_en = reset;
  assign cache_data__T_181_data = 32'h0;
  assign cache_data__T_181_addr = 8'hab;
  assign cache_data__T_181_mask = 1'h0;
  assign cache_data__T_181_en = reset;
  assign cache_data__T_182_data = 32'h0;
  assign cache_data__T_182_addr = 8'hac;
  assign cache_data__T_182_mask = 1'h0;
  assign cache_data__T_182_en = reset;
  assign cache_data__T_183_data = 32'h0;
  assign cache_data__T_183_addr = 8'had;
  assign cache_data__T_183_mask = 1'h0;
  assign cache_data__T_183_en = reset;
  assign cache_data__T_184_data = 32'h0;
  assign cache_data__T_184_addr = 8'hae;
  assign cache_data__T_184_mask = 1'h0;
  assign cache_data__T_184_en = reset;
  assign cache_data__T_185_data = 32'h0;
  assign cache_data__T_185_addr = 8'haf;
  assign cache_data__T_185_mask = 1'h0;
  assign cache_data__T_185_en = reset;
  assign cache_data__T_186_data = 32'h0;
  assign cache_data__T_186_addr = 8'hb0;
  assign cache_data__T_186_mask = 1'h0;
  assign cache_data__T_186_en = reset;
  assign cache_data__T_187_data = 32'h0;
  assign cache_data__T_187_addr = 8'hb1;
  assign cache_data__T_187_mask = 1'h0;
  assign cache_data__T_187_en = reset;
  assign cache_data__T_188_data = 32'h0;
  assign cache_data__T_188_addr = 8'hb2;
  assign cache_data__T_188_mask = 1'h0;
  assign cache_data__T_188_en = reset;
  assign cache_data__T_189_data = 32'h0;
  assign cache_data__T_189_addr = 8'hb3;
  assign cache_data__T_189_mask = 1'h0;
  assign cache_data__T_189_en = reset;
  assign cache_data__T_190_data = 32'h0;
  assign cache_data__T_190_addr = 8'hb4;
  assign cache_data__T_190_mask = 1'h0;
  assign cache_data__T_190_en = reset;
  assign cache_data__T_191_data = 32'h0;
  assign cache_data__T_191_addr = 8'hb5;
  assign cache_data__T_191_mask = 1'h0;
  assign cache_data__T_191_en = reset;
  assign cache_data__T_192_data = 32'h0;
  assign cache_data__T_192_addr = 8'hb6;
  assign cache_data__T_192_mask = 1'h0;
  assign cache_data__T_192_en = reset;
  assign cache_data__T_193_data = 32'h0;
  assign cache_data__T_193_addr = 8'hb7;
  assign cache_data__T_193_mask = 1'h0;
  assign cache_data__T_193_en = reset;
  assign cache_data__T_194_data = 32'h0;
  assign cache_data__T_194_addr = 8'hb8;
  assign cache_data__T_194_mask = 1'h0;
  assign cache_data__T_194_en = reset;
  assign cache_data__T_195_data = 32'h0;
  assign cache_data__T_195_addr = 8'hb9;
  assign cache_data__T_195_mask = 1'h0;
  assign cache_data__T_195_en = reset;
  assign cache_data__T_196_data = 32'h0;
  assign cache_data__T_196_addr = 8'hba;
  assign cache_data__T_196_mask = 1'h0;
  assign cache_data__T_196_en = reset;
  assign cache_data__T_197_data = 32'h0;
  assign cache_data__T_197_addr = 8'hbb;
  assign cache_data__T_197_mask = 1'h0;
  assign cache_data__T_197_en = reset;
  assign cache_data__T_198_data = 32'h0;
  assign cache_data__T_198_addr = 8'hbc;
  assign cache_data__T_198_mask = 1'h0;
  assign cache_data__T_198_en = reset;
  assign cache_data__T_199_data = 32'h0;
  assign cache_data__T_199_addr = 8'hbd;
  assign cache_data__T_199_mask = 1'h0;
  assign cache_data__T_199_en = reset;
  assign cache_data__T_200_data = 32'h0;
  assign cache_data__T_200_addr = 8'hbe;
  assign cache_data__T_200_mask = 1'h0;
  assign cache_data__T_200_en = reset;
  assign cache_data__T_201_data = 32'h0;
  assign cache_data__T_201_addr = 8'hbf;
  assign cache_data__T_201_mask = 1'h0;
  assign cache_data__T_201_en = reset;
  assign cache_data__T_202_data = 32'h0;
  assign cache_data__T_202_addr = 8'hc0;
  assign cache_data__T_202_mask = 1'h0;
  assign cache_data__T_202_en = reset;
  assign cache_data__T_203_data = 32'h0;
  assign cache_data__T_203_addr = 8'hc1;
  assign cache_data__T_203_mask = 1'h0;
  assign cache_data__T_203_en = reset;
  assign cache_data__T_204_data = 32'h0;
  assign cache_data__T_204_addr = 8'hc2;
  assign cache_data__T_204_mask = 1'h0;
  assign cache_data__T_204_en = reset;
  assign cache_data__T_205_data = 32'h0;
  assign cache_data__T_205_addr = 8'hc3;
  assign cache_data__T_205_mask = 1'h0;
  assign cache_data__T_205_en = reset;
  assign cache_data__T_206_data = 32'h0;
  assign cache_data__T_206_addr = 8'hc4;
  assign cache_data__T_206_mask = 1'h0;
  assign cache_data__T_206_en = reset;
  assign cache_data__T_207_data = 32'h0;
  assign cache_data__T_207_addr = 8'hc5;
  assign cache_data__T_207_mask = 1'h0;
  assign cache_data__T_207_en = reset;
  assign cache_data__T_208_data = 32'h0;
  assign cache_data__T_208_addr = 8'hc6;
  assign cache_data__T_208_mask = 1'h0;
  assign cache_data__T_208_en = reset;
  assign cache_data__T_209_data = 32'h0;
  assign cache_data__T_209_addr = 8'hc7;
  assign cache_data__T_209_mask = 1'h0;
  assign cache_data__T_209_en = reset;
  assign cache_data__T_210_data = 32'h0;
  assign cache_data__T_210_addr = 8'hc8;
  assign cache_data__T_210_mask = 1'h0;
  assign cache_data__T_210_en = reset;
  assign cache_data__T_211_data = 32'h0;
  assign cache_data__T_211_addr = 8'hc9;
  assign cache_data__T_211_mask = 1'h0;
  assign cache_data__T_211_en = reset;
  assign cache_data__T_212_data = 32'h0;
  assign cache_data__T_212_addr = 8'hca;
  assign cache_data__T_212_mask = 1'h0;
  assign cache_data__T_212_en = reset;
  assign cache_data__T_213_data = 32'h0;
  assign cache_data__T_213_addr = 8'hcb;
  assign cache_data__T_213_mask = 1'h0;
  assign cache_data__T_213_en = reset;
  assign cache_data__T_214_data = 32'h0;
  assign cache_data__T_214_addr = 8'hcc;
  assign cache_data__T_214_mask = 1'h0;
  assign cache_data__T_214_en = reset;
  assign cache_data__T_215_data = 32'h0;
  assign cache_data__T_215_addr = 8'hcd;
  assign cache_data__T_215_mask = 1'h0;
  assign cache_data__T_215_en = reset;
  assign cache_data__T_216_data = 32'h0;
  assign cache_data__T_216_addr = 8'hce;
  assign cache_data__T_216_mask = 1'h0;
  assign cache_data__T_216_en = reset;
  assign cache_data__T_217_data = 32'h0;
  assign cache_data__T_217_addr = 8'hcf;
  assign cache_data__T_217_mask = 1'h0;
  assign cache_data__T_217_en = reset;
  assign cache_data__T_218_data = 32'h0;
  assign cache_data__T_218_addr = 8'hd0;
  assign cache_data__T_218_mask = 1'h0;
  assign cache_data__T_218_en = reset;
  assign cache_data__T_219_data = 32'h0;
  assign cache_data__T_219_addr = 8'hd1;
  assign cache_data__T_219_mask = 1'h0;
  assign cache_data__T_219_en = reset;
  assign cache_data__T_220_data = 32'h0;
  assign cache_data__T_220_addr = 8'hd2;
  assign cache_data__T_220_mask = 1'h0;
  assign cache_data__T_220_en = reset;
  assign cache_data__T_221_data = 32'h0;
  assign cache_data__T_221_addr = 8'hd3;
  assign cache_data__T_221_mask = 1'h0;
  assign cache_data__T_221_en = reset;
  assign cache_data__T_222_data = 32'h0;
  assign cache_data__T_222_addr = 8'hd4;
  assign cache_data__T_222_mask = 1'h0;
  assign cache_data__T_222_en = reset;
  assign cache_data__T_223_data = 32'h0;
  assign cache_data__T_223_addr = 8'hd5;
  assign cache_data__T_223_mask = 1'h0;
  assign cache_data__T_223_en = reset;
  assign cache_data__T_224_data = 32'h0;
  assign cache_data__T_224_addr = 8'hd6;
  assign cache_data__T_224_mask = 1'h0;
  assign cache_data__T_224_en = reset;
  assign cache_data__T_225_data = 32'h0;
  assign cache_data__T_225_addr = 8'hd7;
  assign cache_data__T_225_mask = 1'h0;
  assign cache_data__T_225_en = reset;
  assign cache_data__T_226_data = 32'h0;
  assign cache_data__T_226_addr = 8'hd8;
  assign cache_data__T_226_mask = 1'h0;
  assign cache_data__T_226_en = reset;
  assign cache_data__T_227_data = 32'h0;
  assign cache_data__T_227_addr = 8'hd9;
  assign cache_data__T_227_mask = 1'h0;
  assign cache_data__T_227_en = reset;
  assign cache_data__T_228_data = 32'h0;
  assign cache_data__T_228_addr = 8'hda;
  assign cache_data__T_228_mask = 1'h0;
  assign cache_data__T_228_en = reset;
  assign cache_data__T_229_data = 32'h0;
  assign cache_data__T_229_addr = 8'hdb;
  assign cache_data__T_229_mask = 1'h0;
  assign cache_data__T_229_en = reset;
  assign cache_data__T_230_data = 32'h0;
  assign cache_data__T_230_addr = 8'hdc;
  assign cache_data__T_230_mask = 1'h0;
  assign cache_data__T_230_en = reset;
  assign cache_data__T_231_data = 32'h0;
  assign cache_data__T_231_addr = 8'hdd;
  assign cache_data__T_231_mask = 1'h0;
  assign cache_data__T_231_en = reset;
  assign cache_data__T_232_data = 32'h0;
  assign cache_data__T_232_addr = 8'hde;
  assign cache_data__T_232_mask = 1'h0;
  assign cache_data__T_232_en = reset;
  assign cache_data__T_233_data = 32'h0;
  assign cache_data__T_233_addr = 8'hdf;
  assign cache_data__T_233_mask = 1'h0;
  assign cache_data__T_233_en = reset;
  assign cache_data__T_234_data = 32'h0;
  assign cache_data__T_234_addr = 8'he0;
  assign cache_data__T_234_mask = 1'h0;
  assign cache_data__T_234_en = reset;
  assign cache_data__T_235_data = 32'h0;
  assign cache_data__T_235_addr = 8'he1;
  assign cache_data__T_235_mask = 1'h0;
  assign cache_data__T_235_en = reset;
  assign cache_data__T_236_data = 32'h0;
  assign cache_data__T_236_addr = 8'he2;
  assign cache_data__T_236_mask = 1'h0;
  assign cache_data__T_236_en = reset;
  assign cache_data__T_237_data = 32'h0;
  assign cache_data__T_237_addr = 8'he3;
  assign cache_data__T_237_mask = 1'h0;
  assign cache_data__T_237_en = reset;
  assign cache_data__T_238_data = 32'h0;
  assign cache_data__T_238_addr = 8'he4;
  assign cache_data__T_238_mask = 1'h0;
  assign cache_data__T_238_en = reset;
  assign cache_data__T_239_data = 32'h0;
  assign cache_data__T_239_addr = 8'he5;
  assign cache_data__T_239_mask = 1'h0;
  assign cache_data__T_239_en = reset;
  assign cache_data__T_240_data = 32'h0;
  assign cache_data__T_240_addr = 8'he6;
  assign cache_data__T_240_mask = 1'h0;
  assign cache_data__T_240_en = reset;
  assign cache_data__T_241_data = 32'h0;
  assign cache_data__T_241_addr = 8'he7;
  assign cache_data__T_241_mask = 1'h0;
  assign cache_data__T_241_en = reset;
  assign cache_data__T_242_data = 32'h0;
  assign cache_data__T_242_addr = 8'he8;
  assign cache_data__T_242_mask = 1'h0;
  assign cache_data__T_242_en = reset;
  assign cache_data__T_243_data = 32'h0;
  assign cache_data__T_243_addr = 8'he9;
  assign cache_data__T_243_mask = 1'h0;
  assign cache_data__T_243_en = reset;
  assign cache_data__T_244_data = 32'h0;
  assign cache_data__T_244_addr = 8'hea;
  assign cache_data__T_244_mask = 1'h0;
  assign cache_data__T_244_en = reset;
  assign cache_data__T_245_data = 32'h0;
  assign cache_data__T_245_addr = 8'heb;
  assign cache_data__T_245_mask = 1'h0;
  assign cache_data__T_245_en = reset;
  assign cache_data__T_246_data = 32'h0;
  assign cache_data__T_246_addr = 8'hec;
  assign cache_data__T_246_mask = 1'h0;
  assign cache_data__T_246_en = reset;
  assign cache_data__T_247_data = 32'h0;
  assign cache_data__T_247_addr = 8'hed;
  assign cache_data__T_247_mask = 1'h0;
  assign cache_data__T_247_en = reset;
  assign cache_data__T_248_data = 32'h0;
  assign cache_data__T_248_addr = 8'hee;
  assign cache_data__T_248_mask = 1'h0;
  assign cache_data__T_248_en = reset;
  assign cache_data__T_249_data = 32'h0;
  assign cache_data__T_249_addr = 8'hef;
  assign cache_data__T_249_mask = 1'h0;
  assign cache_data__T_249_en = reset;
  assign cache_data__T_250_data = 32'h0;
  assign cache_data__T_250_addr = 8'hf0;
  assign cache_data__T_250_mask = 1'h0;
  assign cache_data__T_250_en = reset;
  assign cache_data__T_251_data = 32'h0;
  assign cache_data__T_251_addr = 8'hf1;
  assign cache_data__T_251_mask = 1'h0;
  assign cache_data__T_251_en = reset;
  assign cache_data__T_252_data = 32'h0;
  assign cache_data__T_252_addr = 8'hf2;
  assign cache_data__T_252_mask = 1'h0;
  assign cache_data__T_252_en = reset;
  assign cache_data__T_253_data = 32'h0;
  assign cache_data__T_253_addr = 8'hf3;
  assign cache_data__T_253_mask = 1'h0;
  assign cache_data__T_253_en = reset;
  assign cache_data__T_254_data = 32'h0;
  assign cache_data__T_254_addr = 8'hf4;
  assign cache_data__T_254_mask = 1'h0;
  assign cache_data__T_254_en = reset;
  assign cache_data__T_255_data = 32'h0;
  assign cache_data__T_255_addr = 8'hf5;
  assign cache_data__T_255_mask = 1'h0;
  assign cache_data__T_255_en = reset;
  assign cache_data__T_256_data = 32'h0;
  assign cache_data__T_256_addr = 8'hf6;
  assign cache_data__T_256_mask = 1'h0;
  assign cache_data__T_256_en = reset;
  assign cache_data__T_257_data = 32'h0;
  assign cache_data__T_257_addr = 8'hf7;
  assign cache_data__T_257_mask = 1'h0;
  assign cache_data__T_257_en = reset;
  assign cache_data__T_258_data = 32'h0;
  assign cache_data__T_258_addr = 8'hf8;
  assign cache_data__T_258_mask = 1'h0;
  assign cache_data__T_258_en = reset;
  assign cache_data__T_259_data = 32'h0;
  assign cache_data__T_259_addr = 8'hf9;
  assign cache_data__T_259_mask = 1'h0;
  assign cache_data__T_259_en = reset;
  assign cache_data__T_260_data = 32'h0;
  assign cache_data__T_260_addr = 8'hfa;
  assign cache_data__T_260_mask = 1'h0;
  assign cache_data__T_260_en = reset;
  assign cache_data__T_261_data = 32'h0;
  assign cache_data__T_261_addr = 8'hfb;
  assign cache_data__T_261_mask = 1'h0;
  assign cache_data__T_261_en = reset;
  assign cache_data__T_262_data = 32'h0;
  assign cache_data__T_262_addr = 8'hfc;
  assign cache_data__T_262_mask = 1'h0;
  assign cache_data__T_262_en = reset;
  assign cache_data__T_263_data = 32'h0;
  assign cache_data__T_263_addr = 8'hfd;
  assign cache_data__T_263_mask = 1'h0;
  assign cache_data__T_263_en = reset;
  assign cache_data__T_264_data = 32'h0;
  assign cache_data__T_264_addr = 8'hfe;
  assign cache_data__T_264_mask = 1'h0;
  assign cache_data__T_264_en = reset;
  assign cache_data__T_265_data = 32'h0;
  assign cache_data__T_265_addr = 8'hff;
  assign cache_data__T_265_mask = 1'h0;
  assign cache_data__T_265_en = reset;
  assign cache_data_s1_entry_w_data = io_out_resp_bits_data;
  assign cache_data_s1_entry_w_addr = s1_in_addr[7:0];
  assign cache_data_s1_entry_w_mask = s1_resp & _T_285;
  assign cache_data_s1_entry_w_en = s1_resp & _T_285;
  assign io_in_req_ready = s0_out_ready | _T_268; // @[icache.scala 117:19]
  assign io_in_resp_valid = _T_290 & _T_291; // @[icache.scala 137:20]
  assign io_in_resp_bits_data = cache_data_s1_entry_r_data; // @[icache.scala 138:24]
  assign io_out_req_valid = s1_req; // @[icache.scala 158:20]
  assign io_out_req_bits_is_cached = s1_in_is_cached; // @[icache.scala 159:19]
  assign io_out_req_bits_addr = s1_in_addr; // @[icache.scala 159:19]
  assign io_out_req_bits_len = s1_in_len; // @[icache.scala 159:19]
  assign io_out_req_bits_strb = s1_in_strb; // @[icache.scala 159:19]
  assign io_out_resp_ready = 1'h1; // @[icache.scala 160:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    cache_v[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    cache_tag[initvar] = _RAND_1[23:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    cache_data[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  s0_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  s0_in_is_cached = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  s0_in_addr = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  s0_in_len = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  s0_in_strb = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  s1_in_addr = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  s1_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  s1_in_is_cached = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  s1_in_len = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  s1_in_strb = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  s1_req = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  s1_resp = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  s1_ex_wait = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(cache_v__T_8_en & cache_v__T_8_mask) begin
      cache_v[cache_v__T_8_addr] <= cache_v__T_8_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_10_en & cache_v__T_10_mask) begin
      cache_v[cache_v__T_10_addr] <= cache_v__T_10_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_11_en & cache_v__T_11_mask) begin
      cache_v[cache_v__T_11_addr] <= cache_v__T_11_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_12_en & cache_v__T_12_mask) begin
      cache_v[cache_v__T_12_addr] <= cache_v__T_12_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_13_en & cache_v__T_13_mask) begin
      cache_v[cache_v__T_13_addr] <= cache_v__T_13_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_14_en & cache_v__T_14_mask) begin
      cache_v[cache_v__T_14_addr] <= cache_v__T_14_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_15_en & cache_v__T_15_mask) begin
      cache_v[cache_v__T_15_addr] <= cache_v__T_15_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_16_en & cache_v__T_16_mask) begin
      cache_v[cache_v__T_16_addr] <= cache_v__T_16_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_17_en & cache_v__T_17_mask) begin
      cache_v[cache_v__T_17_addr] <= cache_v__T_17_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_18_en & cache_v__T_18_mask) begin
      cache_v[cache_v__T_18_addr] <= cache_v__T_18_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_19_en & cache_v__T_19_mask) begin
      cache_v[cache_v__T_19_addr] <= cache_v__T_19_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_20_en & cache_v__T_20_mask) begin
      cache_v[cache_v__T_20_addr] <= cache_v__T_20_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_21_en & cache_v__T_21_mask) begin
      cache_v[cache_v__T_21_addr] <= cache_v__T_21_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_22_en & cache_v__T_22_mask) begin
      cache_v[cache_v__T_22_addr] <= cache_v__T_22_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_23_en & cache_v__T_23_mask) begin
      cache_v[cache_v__T_23_addr] <= cache_v__T_23_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_24_en & cache_v__T_24_mask) begin
      cache_v[cache_v__T_24_addr] <= cache_v__T_24_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_25_en & cache_v__T_25_mask) begin
      cache_v[cache_v__T_25_addr] <= cache_v__T_25_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_26_en & cache_v__T_26_mask) begin
      cache_v[cache_v__T_26_addr] <= cache_v__T_26_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_27_en & cache_v__T_27_mask) begin
      cache_v[cache_v__T_27_addr] <= cache_v__T_27_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_28_en & cache_v__T_28_mask) begin
      cache_v[cache_v__T_28_addr] <= cache_v__T_28_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_29_en & cache_v__T_29_mask) begin
      cache_v[cache_v__T_29_addr] <= cache_v__T_29_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_30_en & cache_v__T_30_mask) begin
      cache_v[cache_v__T_30_addr] <= cache_v__T_30_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_31_en & cache_v__T_31_mask) begin
      cache_v[cache_v__T_31_addr] <= cache_v__T_31_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_32_en & cache_v__T_32_mask) begin
      cache_v[cache_v__T_32_addr] <= cache_v__T_32_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_33_en & cache_v__T_33_mask) begin
      cache_v[cache_v__T_33_addr] <= cache_v__T_33_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_34_en & cache_v__T_34_mask) begin
      cache_v[cache_v__T_34_addr] <= cache_v__T_34_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_35_en & cache_v__T_35_mask) begin
      cache_v[cache_v__T_35_addr] <= cache_v__T_35_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_36_en & cache_v__T_36_mask) begin
      cache_v[cache_v__T_36_addr] <= cache_v__T_36_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_37_en & cache_v__T_37_mask) begin
      cache_v[cache_v__T_37_addr] <= cache_v__T_37_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_38_en & cache_v__T_38_mask) begin
      cache_v[cache_v__T_38_addr] <= cache_v__T_38_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_39_en & cache_v__T_39_mask) begin
      cache_v[cache_v__T_39_addr] <= cache_v__T_39_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_40_en & cache_v__T_40_mask) begin
      cache_v[cache_v__T_40_addr] <= cache_v__T_40_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_41_en & cache_v__T_41_mask) begin
      cache_v[cache_v__T_41_addr] <= cache_v__T_41_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_42_en & cache_v__T_42_mask) begin
      cache_v[cache_v__T_42_addr] <= cache_v__T_42_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_43_en & cache_v__T_43_mask) begin
      cache_v[cache_v__T_43_addr] <= cache_v__T_43_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_44_en & cache_v__T_44_mask) begin
      cache_v[cache_v__T_44_addr] <= cache_v__T_44_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_45_en & cache_v__T_45_mask) begin
      cache_v[cache_v__T_45_addr] <= cache_v__T_45_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_46_en & cache_v__T_46_mask) begin
      cache_v[cache_v__T_46_addr] <= cache_v__T_46_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_47_en & cache_v__T_47_mask) begin
      cache_v[cache_v__T_47_addr] <= cache_v__T_47_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_48_en & cache_v__T_48_mask) begin
      cache_v[cache_v__T_48_addr] <= cache_v__T_48_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_49_en & cache_v__T_49_mask) begin
      cache_v[cache_v__T_49_addr] <= cache_v__T_49_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_50_en & cache_v__T_50_mask) begin
      cache_v[cache_v__T_50_addr] <= cache_v__T_50_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_51_en & cache_v__T_51_mask) begin
      cache_v[cache_v__T_51_addr] <= cache_v__T_51_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_52_en & cache_v__T_52_mask) begin
      cache_v[cache_v__T_52_addr] <= cache_v__T_52_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_53_en & cache_v__T_53_mask) begin
      cache_v[cache_v__T_53_addr] <= cache_v__T_53_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_54_en & cache_v__T_54_mask) begin
      cache_v[cache_v__T_54_addr] <= cache_v__T_54_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_55_en & cache_v__T_55_mask) begin
      cache_v[cache_v__T_55_addr] <= cache_v__T_55_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_56_en & cache_v__T_56_mask) begin
      cache_v[cache_v__T_56_addr] <= cache_v__T_56_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_57_en & cache_v__T_57_mask) begin
      cache_v[cache_v__T_57_addr] <= cache_v__T_57_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_58_en & cache_v__T_58_mask) begin
      cache_v[cache_v__T_58_addr] <= cache_v__T_58_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_59_en & cache_v__T_59_mask) begin
      cache_v[cache_v__T_59_addr] <= cache_v__T_59_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_60_en & cache_v__T_60_mask) begin
      cache_v[cache_v__T_60_addr] <= cache_v__T_60_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_61_en & cache_v__T_61_mask) begin
      cache_v[cache_v__T_61_addr] <= cache_v__T_61_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_62_en & cache_v__T_62_mask) begin
      cache_v[cache_v__T_62_addr] <= cache_v__T_62_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_63_en & cache_v__T_63_mask) begin
      cache_v[cache_v__T_63_addr] <= cache_v__T_63_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_64_en & cache_v__T_64_mask) begin
      cache_v[cache_v__T_64_addr] <= cache_v__T_64_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_65_en & cache_v__T_65_mask) begin
      cache_v[cache_v__T_65_addr] <= cache_v__T_65_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_66_en & cache_v__T_66_mask) begin
      cache_v[cache_v__T_66_addr] <= cache_v__T_66_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_67_en & cache_v__T_67_mask) begin
      cache_v[cache_v__T_67_addr] <= cache_v__T_67_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_68_en & cache_v__T_68_mask) begin
      cache_v[cache_v__T_68_addr] <= cache_v__T_68_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_69_en & cache_v__T_69_mask) begin
      cache_v[cache_v__T_69_addr] <= cache_v__T_69_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_70_en & cache_v__T_70_mask) begin
      cache_v[cache_v__T_70_addr] <= cache_v__T_70_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_71_en & cache_v__T_71_mask) begin
      cache_v[cache_v__T_71_addr] <= cache_v__T_71_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_72_en & cache_v__T_72_mask) begin
      cache_v[cache_v__T_72_addr] <= cache_v__T_72_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_73_en & cache_v__T_73_mask) begin
      cache_v[cache_v__T_73_addr] <= cache_v__T_73_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_74_en & cache_v__T_74_mask) begin
      cache_v[cache_v__T_74_addr] <= cache_v__T_74_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_75_en & cache_v__T_75_mask) begin
      cache_v[cache_v__T_75_addr] <= cache_v__T_75_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_76_en & cache_v__T_76_mask) begin
      cache_v[cache_v__T_76_addr] <= cache_v__T_76_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_77_en & cache_v__T_77_mask) begin
      cache_v[cache_v__T_77_addr] <= cache_v__T_77_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_78_en & cache_v__T_78_mask) begin
      cache_v[cache_v__T_78_addr] <= cache_v__T_78_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_79_en & cache_v__T_79_mask) begin
      cache_v[cache_v__T_79_addr] <= cache_v__T_79_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_80_en & cache_v__T_80_mask) begin
      cache_v[cache_v__T_80_addr] <= cache_v__T_80_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_81_en & cache_v__T_81_mask) begin
      cache_v[cache_v__T_81_addr] <= cache_v__T_81_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_82_en & cache_v__T_82_mask) begin
      cache_v[cache_v__T_82_addr] <= cache_v__T_82_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_83_en & cache_v__T_83_mask) begin
      cache_v[cache_v__T_83_addr] <= cache_v__T_83_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_84_en & cache_v__T_84_mask) begin
      cache_v[cache_v__T_84_addr] <= cache_v__T_84_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_85_en & cache_v__T_85_mask) begin
      cache_v[cache_v__T_85_addr] <= cache_v__T_85_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_86_en & cache_v__T_86_mask) begin
      cache_v[cache_v__T_86_addr] <= cache_v__T_86_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_87_en & cache_v__T_87_mask) begin
      cache_v[cache_v__T_87_addr] <= cache_v__T_87_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_88_en & cache_v__T_88_mask) begin
      cache_v[cache_v__T_88_addr] <= cache_v__T_88_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_89_en & cache_v__T_89_mask) begin
      cache_v[cache_v__T_89_addr] <= cache_v__T_89_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_90_en & cache_v__T_90_mask) begin
      cache_v[cache_v__T_90_addr] <= cache_v__T_90_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_91_en & cache_v__T_91_mask) begin
      cache_v[cache_v__T_91_addr] <= cache_v__T_91_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_92_en & cache_v__T_92_mask) begin
      cache_v[cache_v__T_92_addr] <= cache_v__T_92_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_93_en & cache_v__T_93_mask) begin
      cache_v[cache_v__T_93_addr] <= cache_v__T_93_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_94_en & cache_v__T_94_mask) begin
      cache_v[cache_v__T_94_addr] <= cache_v__T_94_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_95_en & cache_v__T_95_mask) begin
      cache_v[cache_v__T_95_addr] <= cache_v__T_95_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_96_en & cache_v__T_96_mask) begin
      cache_v[cache_v__T_96_addr] <= cache_v__T_96_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_97_en & cache_v__T_97_mask) begin
      cache_v[cache_v__T_97_addr] <= cache_v__T_97_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_98_en & cache_v__T_98_mask) begin
      cache_v[cache_v__T_98_addr] <= cache_v__T_98_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_99_en & cache_v__T_99_mask) begin
      cache_v[cache_v__T_99_addr] <= cache_v__T_99_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_100_en & cache_v__T_100_mask) begin
      cache_v[cache_v__T_100_addr] <= cache_v__T_100_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_101_en & cache_v__T_101_mask) begin
      cache_v[cache_v__T_101_addr] <= cache_v__T_101_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_102_en & cache_v__T_102_mask) begin
      cache_v[cache_v__T_102_addr] <= cache_v__T_102_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_103_en & cache_v__T_103_mask) begin
      cache_v[cache_v__T_103_addr] <= cache_v__T_103_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_104_en & cache_v__T_104_mask) begin
      cache_v[cache_v__T_104_addr] <= cache_v__T_104_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_105_en & cache_v__T_105_mask) begin
      cache_v[cache_v__T_105_addr] <= cache_v__T_105_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_106_en & cache_v__T_106_mask) begin
      cache_v[cache_v__T_106_addr] <= cache_v__T_106_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_107_en & cache_v__T_107_mask) begin
      cache_v[cache_v__T_107_addr] <= cache_v__T_107_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_108_en & cache_v__T_108_mask) begin
      cache_v[cache_v__T_108_addr] <= cache_v__T_108_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_109_en & cache_v__T_109_mask) begin
      cache_v[cache_v__T_109_addr] <= cache_v__T_109_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_110_en & cache_v__T_110_mask) begin
      cache_v[cache_v__T_110_addr] <= cache_v__T_110_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_111_en & cache_v__T_111_mask) begin
      cache_v[cache_v__T_111_addr] <= cache_v__T_111_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_112_en & cache_v__T_112_mask) begin
      cache_v[cache_v__T_112_addr] <= cache_v__T_112_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_113_en & cache_v__T_113_mask) begin
      cache_v[cache_v__T_113_addr] <= cache_v__T_113_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_114_en & cache_v__T_114_mask) begin
      cache_v[cache_v__T_114_addr] <= cache_v__T_114_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_115_en & cache_v__T_115_mask) begin
      cache_v[cache_v__T_115_addr] <= cache_v__T_115_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_116_en & cache_v__T_116_mask) begin
      cache_v[cache_v__T_116_addr] <= cache_v__T_116_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_117_en & cache_v__T_117_mask) begin
      cache_v[cache_v__T_117_addr] <= cache_v__T_117_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_118_en & cache_v__T_118_mask) begin
      cache_v[cache_v__T_118_addr] <= cache_v__T_118_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_119_en & cache_v__T_119_mask) begin
      cache_v[cache_v__T_119_addr] <= cache_v__T_119_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_120_en & cache_v__T_120_mask) begin
      cache_v[cache_v__T_120_addr] <= cache_v__T_120_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_121_en & cache_v__T_121_mask) begin
      cache_v[cache_v__T_121_addr] <= cache_v__T_121_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_122_en & cache_v__T_122_mask) begin
      cache_v[cache_v__T_122_addr] <= cache_v__T_122_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_123_en & cache_v__T_123_mask) begin
      cache_v[cache_v__T_123_addr] <= cache_v__T_123_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_124_en & cache_v__T_124_mask) begin
      cache_v[cache_v__T_124_addr] <= cache_v__T_124_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_125_en & cache_v__T_125_mask) begin
      cache_v[cache_v__T_125_addr] <= cache_v__T_125_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_126_en & cache_v__T_126_mask) begin
      cache_v[cache_v__T_126_addr] <= cache_v__T_126_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_127_en & cache_v__T_127_mask) begin
      cache_v[cache_v__T_127_addr] <= cache_v__T_127_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_128_en & cache_v__T_128_mask) begin
      cache_v[cache_v__T_128_addr] <= cache_v__T_128_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_129_en & cache_v__T_129_mask) begin
      cache_v[cache_v__T_129_addr] <= cache_v__T_129_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_130_en & cache_v__T_130_mask) begin
      cache_v[cache_v__T_130_addr] <= cache_v__T_130_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_131_en & cache_v__T_131_mask) begin
      cache_v[cache_v__T_131_addr] <= cache_v__T_131_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_132_en & cache_v__T_132_mask) begin
      cache_v[cache_v__T_132_addr] <= cache_v__T_132_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_133_en & cache_v__T_133_mask) begin
      cache_v[cache_v__T_133_addr] <= cache_v__T_133_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_134_en & cache_v__T_134_mask) begin
      cache_v[cache_v__T_134_addr] <= cache_v__T_134_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_135_en & cache_v__T_135_mask) begin
      cache_v[cache_v__T_135_addr] <= cache_v__T_135_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_136_en & cache_v__T_136_mask) begin
      cache_v[cache_v__T_136_addr] <= cache_v__T_136_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_137_en & cache_v__T_137_mask) begin
      cache_v[cache_v__T_137_addr] <= cache_v__T_137_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_138_en & cache_v__T_138_mask) begin
      cache_v[cache_v__T_138_addr] <= cache_v__T_138_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_139_en & cache_v__T_139_mask) begin
      cache_v[cache_v__T_139_addr] <= cache_v__T_139_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_140_en & cache_v__T_140_mask) begin
      cache_v[cache_v__T_140_addr] <= cache_v__T_140_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_141_en & cache_v__T_141_mask) begin
      cache_v[cache_v__T_141_addr] <= cache_v__T_141_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_142_en & cache_v__T_142_mask) begin
      cache_v[cache_v__T_142_addr] <= cache_v__T_142_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_143_en & cache_v__T_143_mask) begin
      cache_v[cache_v__T_143_addr] <= cache_v__T_143_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_144_en & cache_v__T_144_mask) begin
      cache_v[cache_v__T_144_addr] <= cache_v__T_144_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_145_en & cache_v__T_145_mask) begin
      cache_v[cache_v__T_145_addr] <= cache_v__T_145_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_146_en & cache_v__T_146_mask) begin
      cache_v[cache_v__T_146_addr] <= cache_v__T_146_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_147_en & cache_v__T_147_mask) begin
      cache_v[cache_v__T_147_addr] <= cache_v__T_147_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_148_en & cache_v__T_148_mask) begin
      cache_v[cache_v__T_148_addr] <= cache_v__T_148_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_149_en & cache_v__T_149_mask) begin
      cache_v[cache_v__T_149_addr] <= cache_v__T_149_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_150_en & cache_v__T_150_mask) begin
      cache_v[cache_v__T_150_addr] <= cache_v__T_150_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_151_en & cache_v__T_151_mask) begin
      cache_v[cache_v__T_151_addr] <= cache_v__T_151_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_152_en & cache_v__T_152_mask) begin
      cache_v[cache_v__T_152_addr] <= cache_v__T_152_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_153_en & cache_v__T_153_mask) begin
      cache_v[cache_v__T_153_addr] <= cache_v__T_153_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_154_en & cache_v__T_154_mask) begin
      cache_v[cache_v__T_154_addr] <= cache_v__T_154_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_155_en & cache_v__T_155_mask) begin
      cache_v[cache_v__T_155_addr] <= cache_v__T_155_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_156_en & cache_v__T_156_mask) begin
      cache_v[cache_v__T_156_addr] <= cache_v__T_156_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_157_en & cache_v__T_157_mask) begin
      cache_v[cache_v__T_157_addr] <= cache_v__T_157_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_158_en & cache_v__T_158_mask) begin
      cache_v[cache_v__T_158_addr] <= cache_v__T_158_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_159_en & cache_v__T_159_mask) begin
      cache_v[cache_v__T_159_addr] <= cache_v__T_159_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_160_en & cache_v__T_160_mask) begin
      cache_v[cache_v__T_160_addr] <= cache_v__T_160_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_161_en & cache_v__T_161_mask) begin
      cache_v[cache_v__T_161_addr] <= cache_v__T_161_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_162_en & cache_v__T_162_mask) begin
      cache_v[cache_v__T_162_addr] <= cache_v__T_162_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_163_en & cache_v__T_163_mask) begin
      cache_v[cache_v__T_163_addr] <= cache_v__T_163_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_164_en & cache_v__T_164_mask) begin
      cache_v[cache_v__T_164_addr] <= cache_v__T_164_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_165_en & cache_v__T_165_mask) begin
      cache_v[cache_v__T_165_addr] <= cache_v__T_165_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_166_en & cache_v__T_166_mask) begin
      cache_v[cache_v__T_166_addr] <= cache_v__T_166_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_167_en & cache_v__T_167_mask) begin
      cache_v[cache_v__T_167_addr] <= cache_v__T_167_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_168_en & cache_v__T_168_mask) begin
      cache_v[cache_v__T_168_addr] <= cache_v__T_168_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_169_en & cache_v__T_169_mask) begin
      cache_v[cache_v__T_169_addr] <= cache_v__T_169_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_170_en & cache_v__T_170_mask) begin
      cache_v[cache_v__T_170_addr] <= cache_v__T_170_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_171_en & cache_v__T_171_mask) begin
      cache_v[cache_v__T_171_addr] <= cache_v__T_171_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_172_en & cache_v__T_172_mask) begin
      cache_v[cache_v__T_172_addr] <= cache_v__T_172_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_173_en & cache_v__T_173_mask) begin
      cache_v[cache_v__T_173_addr] <= cache_v__T_173_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_174_en & cache_v__T_174_mask) begin
      cache_v[cache_v__T_174_addr] <= cache_v__T_174_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_175_en & cache_v__T_175_mask) begin
      cache_v[cache_v__T_175_addr] <= cache_v__T_175_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_176_en & cache_v__T_176_mask) begin
      cache_v[cache_v__T_176_addr] <= cache_v__T_176_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_177_en & cache_v__T_177_mask) begin
      cache_v[cache_v__T_177_addr] <= cache_v__T_177_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_178_en & cache_v__T_178_mask) begin
      cache_v[cache_v__T_178_addr] <= cache_v__T_178_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_179_en & cache_v__T_179_mask) begin
      cache_v[cache_v__T_179_addr] <= cache_v__T_179_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_180_en & cache_v__T_180_mask) begin
      cache_v[cache_v__T_180_addr] <= cache_v__T_180_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_181_en & cache_v__T_181_mask) begin
      cache_v[cache_v__T_181_addr] <= cache_v__T_181_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_182_en & cache_v__T_182_mask) begin
      cache_v[cache_v__T_182_addr] <= cache_v__T_182_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_183_en & cache_v__T_183_mask) begin
      cache_v[cache_v__T_183_addr] <= cache_v__T_183_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_184_en & cache_v__T_184_mask) begin
      cache_v[cache_v__T_184_addr] <= cache_v__T_184_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_185_en & cache_v__T_185_mask) begin
      cache_v[cache_v__T_185_addr] <= cache_v__T_185_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_186_en & cache_v__T_186_mask) begin
      cache_v[cache_v__T_186_addr] <= cache_v__T_186_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_187_en & cache_v__T_187_mask) begin
      cache_v[cache_v__T_187_addr] <= cache_v__T_187_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_188_en & cache_v__T_188_mask) begin
      cache_v[cache_v__T_188_addr] <= cache_v__T_188_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_189_en & cache_v__T_189_mask) begin
      cache_v[cache_v__T_189_addr] <= cache_v__T_189_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_190_en & cache_v__T_190_mask) begin
      cache_v[cache_v__T_190_addr] <= cache_v__T_190_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_191_en & cache_v__T_191_mask) begin
      cache_v[cache_v__T_191_addr] <= cache_v__T_191_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_192_en & cache_v__T_192_mask) begin
      cache_v[cache_v__T_192_addr] <= cache_v__T_192_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_193_en & cache_v__T_193_mask) begin
      cache_v[cache_v__T_193_addr] <= cache_v__T_193_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_194_en & cache_v__T_194_mask) begin
      cache_v[cache_v__T_194_addr] <= cache_v__T_194_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_195_en & cache_v__T_195_mask) begin
      cache_v[cache_v__T_195_addr] <= cache_v__T_195_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_196_en & cache_v__T_196_mask) begin
      cache_v[cache_v__T_196_addr] <= cache_v__T_196_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_197_en & cache_v__T_197_mask) begin
      cache_v[cache_v__T_197_addr] <= cache_v__T_197_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_198_en & cache_v__T_198_mask) begin
      cache_v[cache_v__T_198_addr] <= cache_v__T_198_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_199_en & cache_v__T_199_mask) begin
      cache_v[cache_v__T_199_addr] <= cache_v__T_199_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_200_en & cache_v__T_200_mask) begin
      cache_v[cache_v__T_200_addr] <= cache_v__T_200_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_201_en & cache_v__T_201_mask) begin
      cache_v[cache_v__T_201_addr] <= cache_v__T_201_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_202_en & cache_v__T_202_mask) begin
      cache_v[cache_v__T_202_addr] <= cache_v__T_202_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_203_en & cache_v__T_203_mask) begin
      cache_v[cache_v__T_203_addr] <= cache_v__T_203_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_204_en & cache_v__T_204_mask) begin
      cache_v[cache_v__T_204_addr] <= cache_v__T_204_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_205_en & cache_v__T_205_mask) begin
      cache_v[cache_v__T_205_addr] <= cache_v__T_205_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_206_en & cache_v__T_206_mask) begin
      cache_v[cache_v__T_206_addr] <= cache_v__T_206_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_207_en & cache_v__T_207_mask) begin
      cache_v[cache_v__T_207_addr] <= cache_v__T_207_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_208_en & cache_v__T_208_mask) begin
      cache_v[cache_v__T_208_addr] <= cache_v__T_208_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_209_en & cache_v__T_209_mask) begin
      cache_v[cache_v__T_209_addr] <= cache_v__T_209_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_210_en & cache_v__T_210_mask) begin
      cache_v[cache_v__T_210_addr] <= cache_v__T_210_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_211_en & cache_v__T_211_mask) begin
      cache_v[cache_v__T_211_addr] <= cache_v__T_211_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_212_en & cache_v__T_212_mask) begin
      cache_v[cache_v__T_212_addr] <= cache_v__T_212_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_213_en & cache_v__T_213_mask) begin
      cache_v[cache_v__T_213_addr] <= cache_v__T_213_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_214_en & cache_v__T_214_mask) begin
      cache_v[cache_v__T_214_addr] <= cache_v__T_214_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_215_en & cache_v__T_215_mask) begin
      cache_v[cache_v__T_215_addr] <= cache_v__T_215_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_216_en & cache_v__T_216_mask) begin
      cache_v[cache_v__T_216_addr] <= cache_v__T_216_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_217_en & cache_v__T_217_mask) begin
      cache_v[cache_v__T_217_addr] <= cache_v__T_217_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_218_en & cache_v__T_218_mask) begin
      cache_v[cache_v__T_218_addr] <= cache_v__T_218_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_219_en & cache_v__T_219_mask) begin
      cache_v[cache_v__T_219_addr] <= cache_v__T_219_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_220_en & cache_v__T_220_mask) begin
      cache_v[cache_v__T_220_addr] <= cache_v__T_220_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_221_en & cache_v__T_221_mask) begin
      cache_v[cache_v__T_221_addr] <= cache_v__T_221_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_222_en & cache_v__T_222_mask) begin
      cache_v[cache_v__T_222_addr] <= cache_v__T_222_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_223_en & cache_v__T_223_mask) begin
      cache_v[cache_v__T_223_addr] <= cache_v__T_223_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_224_en & cache_v__T_224_mask) begin
      cache_v[cache_v__T_224_addr] <= cache_v__T_224_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_225_en & cache_v__T_225_mask) begin
      cache_v[cache_v__T_225_addr] <= cache_v__T_225_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_226_en & cache_v__T_226_mask) begin
      cache_v[cache_v__T_226_addr] <= cache_v__T_226_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_227_en & cache_v__T_227_mask) begin
      cache_v[cache_v__T_227_addr] <= cache_v__T_227_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_228_en & cache_v__T_228_mask) begin
      cache_v[cache_v__T_228_addr] <= cache_v__T_228_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_229_en & cache_v__T_229_mask) begin
      cache_v[cache_v__T_229_addr] <= cache_v__T_229_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_230_en & cache_v__T_230_mask) begin
      cache_v[cache_v__T_230_addr] <= cache_v__T_230_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_231_en & cache_v__T_231_mask) begin
      cache_v[cache_v__T_231_addr] <= cache_v__T_231_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_232_en & cache_v__T_232_mask) begin
      cache_v[cache_v__T_232_addr] <= cache_v__T_232_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_233_en & cache_v__T_233_mask) begin
      cache_v[cache_v__T_233_addr] <= cache_v__T_233_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_234_en & cache_v__T_234_mask) begin
      cache_v[cache_v__T_234_addr] <= cache_v__T_234_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_235_en & cache_v__T_235_mask) begin
      cache_v[cache_v__T_235_addr] <= cache_v__T_235_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_236_en & cache_v__T_236_mask) begin
      cache_v[cache_v__T_236_addr] <= cache_v__T_236_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_237_en & cache_v__T_237_mask) begin
      cache_v[cache_v__T_237_addr] <= cache_v__T_237_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_238_en & cache_v__T_238_mask) begin
      cache_v[cache_v__T_238_addr] <= cache_v__T_238_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_239_en & cache_v__T_239_mask) begin
      cache_v[cache_v__T_239_addr] <= cache_v__T_239_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_240_en & cache_v__T_240_mask) begin
      cache_v[cache_v__T_240_addr] <= cache_v__T_240_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_241_en & cache_v__T_241_mask) begin
      cache_v[cache_v__T_241_addr] <= cache_v__T_241_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_242_en & cache_v__T_242_mask) begin
      cache_v[cache_v__T_242_addr] <= cache_v__T_242_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_243_en & cache_v__T_243_mask) begin
      cache_v[cache_v__T_243_addr] <= cache_v__T_243_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_244_en & cache_v__T_244_mask) begin
      cache_v[cache_v__T_244_addr] <= cache_v__T_244_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_245_en & cache_v__T_245_mask) begin
      cache_v[cache_v__T_245_addr] <= cache_v__T_245_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_246_en & cache_v__T_246_mask) begin
      cache_v[cache_v__T_246_addr] <= cache_v__T_246_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_247_en & cache_v__T_247_mask) begin
      cache_v[cache_v__T_247_addr] <= cache_v__T_247_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_248_en & cache_v__T_248_mask) begin
      cache_v[cache_v__T_248_addr] <= cache_v__T_248_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_249_en & cache_v__T_249_mask) begin
      cache_v[cache_v__T_249_addr] <= cache_v__T_249_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_250_en & cache_v__T_250_mask) begin
      cache_v[cache_v__T_250_addr] <= cache_v__T_250_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_251_en & cache_v__T_251_mask) begin
      cache_v[cache_v__T_251_addr] <= cache_v__T_251_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_252_en & cache_v__T_252_mask) begin
      cache_v[cache_v__T_252_addr] <= cache_v__T_252_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_253_en & cache_v__T_253_mask) begin
      cache_v[cache_v__T_253_addr] <= cache_v__T_253_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_254_en & cache_v__T_254_mask) begin
      cache_v[cache_v__T_254_addr] <= cache_v__T_254_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_255_en & cache_v__T_255_mask) begin
      cache_v[cache_v__T_255_addr] <= cache_v__T_255_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_256_en & cache_v__T_256_mask) begin
      cache_v[cache_v__T_256_addr] <= cache_v__T_256_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_257_en & cache_v__T_257_mask) begin
      cache_v[cache_v__T_257_addr] <= cache_v__T_257_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_258_en & cache_v__T_258_mask) begin
      cache_v[cache_v__T_258_addr] <= cache_v__T_258_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_259_en & cache_v__T_259_mask) begin
      cache_v[cache_v__T_259_addr] <= cache_v__T_259_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_260_en & cache_v__T_260_mask) begin
      cache_v[cache_v__T_260_addr] <= cache_v__T_260_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_261_en & cache_v__T_261_mask) begin
      cache_v[cache_v__T_261_addr] <= cache_v__T_261_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_262_en & cache_v__T_262_mask) begin
      cache_v[cache_v__T_262_addr] <= cache_v__T_262_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_263_en & cache_v__T_263_mask) begin
      cache_v[cache_v__T_263_addr] <= cache_v__T_263_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_264_en & cache_v__T_264_mask) begin
      cache_v[cache_v__T_264_addr] <= cache_v__T_264_data; // @[icache.scala 91:18]
    end
    if(cache_v__T_265_en & cache_v__T_265_mask) begin
      cache_v[cache_v__T_265_addr] <= cache_v__T_265_data; // @[icache.scala 91:18]
    end
    if(cache_v_s1_entry_w_en & cache_v_s1_entry_w_mask) begin
      cache_v[cache_v_s1_entry_w_addr] <= cache_v_s1_entry_w_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_8_en & cache_tag__T_8_mask) begin
      cache_tag[cache_tag__T_8_addr] <= cache_tag__T_8_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_10_en & cache_tag__T_10_mask) begin
      cache_tag[cache_tag__T_10_addr] <= cache_tag__T_10_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_11_en & cache_tag__T_11_mask) begin
      cache_tag[cache_tag__T_11_addr] <= cache_tag__T_11_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_12_en & cache_tag__T_12_mask) begin
      cache_tag[cache_tag__T_12_addr] <= cache_tag__T_12_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_13_en & cache_tag__T_13_mask) begin
      cache_tag[cache_tag__T_13_addr] <= cache_tag__T_13_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_14_en & cache_tag__T_14_mask) begin
      cache_tag[cache_tag__T_14_addr] <= cache_tag__T_14_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_15_en & cache_tag__T_15_mask) begin
      cache_tag[cache_tag__T_15_addr] <= cache_tag__T_15_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_16_en & cache_tag__T_16_mask) begin
      cache_tag[cache_tag__T_16_addr] <= cache_tag__T_16_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_17_en & cache_tag__T_17_mask) begin
      cache_tag[cache_tag__T_17_addr] <= cache_tag__T_17_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_18_en & cache_tag__T_18_mask) begin
      cache_tag[cache_tag__T_18_addr] <= cache_tag__T_18_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_19_en & cache_tag__T_19_mask) begin
      cache_tag[cache_tag__T_19_addr] <= cache_tag__T_19_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_20_en & cache_tag__T_20_mask) begin
      cache_tag[cache_tag__T_20_addr] <= cache_tag__T_20_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_21_en & cache_tag__T_21_mask) begin
      cache_tag[cache_tag__T_21_addr] <= cache_tag__T_21_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_22_en & cache_tag__T_22_mask) begin
      cache_tag[cache_tag__T_22_addr] <= cache_tag__T_22_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_23_en & cache_tag__T_23_mask) begin
      cache_tag[cache_tag__T_23_addr] <= cache_tag__T_23_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_24_en & cache_tag__T_24_mask) begin
      cache_tag[cache_tag__T_24_addr] <= cache_tag__T_24_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_25_en & cache_tag__T_25_mask) begin
      cache_tag[cache_tag__T_25_addr] <= cache_tag__T_25_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_26_en & cache_tag__T_26_mask) begin
      cache_tag[cache_tag__T_26_addr] <= cache_tag__T_26_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_27_en & cache_tag__T_27_mask) begin
      cache_tag[cache_tag__T_27_addr] <= cache_tag__T_27_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_28_en & cache_tag__T_28_mask) begin
      cache_tag[cache_tag__T_28_addr] <= cache_tag__T_28_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_29_en & cache_tag__T_29_mask) begin
      cache_tag[cache_tag__T_29_addr] <= cache_tag__T_29_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_30_en & cache_tag__T_30_mask) begin
      cache_tag[cache_tag__T_30_addr] <= cache_tag__T_30_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_31_en & cache_tag__T_31_mask) begin
      cache_tag[cache_tag__T_31_addr] <= cache_tag__T_31_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_32_en & cache_tag__T_32_mask) begin
      cache_tag[cache_tag__T_32_addr] <= cache_tag__T_32_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_33_en & cache_tag__T_33_mask) begin
      cache_tag[cache_tag__T_33_addr] <= cache_tag__T_33_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_34_en & cache_tag__T_34_mask) begin
      cache_tag[cache_tag__T_34_addr] <= cache_tag__T_34_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_35_en & cache_tag__T_35_mask) begin
      cache_tag[cache_tag__T_35_addr] <= cache_tag__T_35_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_36_en & cache_tag__T_36_mask) begin
      cache_tag[cache_tag__T_36_addr] <= cache_tag__T_36_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_37_en & cache_tag__T_37_mask) begin
      cache_tag[cache_tag__T_37_addr] <= cache_tag__T_37_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_38_en & cache_tag__T_38_mask) begin
      cache_tag[cache_tag__T_38_addr] <= cache_tag__T_38_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_39_en & cache_tag__T_39_mask) begin
      cache_tag[cache_tag__T_39_addr] <= cache_tag__T_39_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_40_en & cache_tag__T_40_mask) begin
      cache_tag[cache_tag__T_40_addr] <= cache_tag__T_40_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_41_en & cache_tag__T_41_mask) begin
      cache_tag[cache_tag__T_41_addr] <= cache_tag__T_41_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_42_en & cache_tag__T_42_mask) begin
      cache_tag[cache_tag__T_42_addr] <= cache_tag__T_42_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_43_en & cache_tag__T_43_mask) begin
      cache_tag[cache_tag__T_43_addr] <= cache_tag__T_43_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_44_en & cache_tag__T_44_mask) begin
      cache_tag[cache_tag__T_44_addr] <= cache_tag__T_44_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_45_en & cache_tag__T_45_mask) begin
      cache_tag[cache_tag__T_45_addr] <= cache_tag__T_45_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_46_en & cache_tag__T_46_mask) begin
      cache_tag[cache_tag__T_46_addr] <= cache_tag__T_46_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_47_en & cache_tag__T_47_mask) begin
      cache_tag[cache_tag__T_47_addr] <= cache_tag__T_47_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_48_en & cache_tag__T_48_mask) begin
      cache_tag[cache_tag__T_48_addr] <= cache_tag__T_48_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_49_en & cache_tag__T_49_mask) begin
      cache_tag[cache_tag__T_49_addr] <= cache_tag__T_49_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_50_en & cache_tag__T_50_mask) begin
      cache_tag[cache_tag__T_50_addr] <= cache_tag__T_50_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_51_en & cache_tag__T_51_mask) begin
      cache_tag[cache_tag__T_51_addr] <= cache_tag__T_51_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_52_en & cache_tag__T_52_mask) begin
      cache_tag[cache_tag__T_52_addr] <= cache_tag__T_52_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_53_en & cache_tag__T_53_mask) begin
      cache_tag[cache_tag__T_53_addr] <= cache_tag__T_53_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_54_en & cache_tag__T_54_mask) begin
      cache_tag[cache_tag__T_54_addr] <= cache_tag__T_54_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_55_en & cache_tag__T_55_mask) begin
      cache_tag[cache_tag__T_55_addr] <= cache_tag__T_55_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_56_en & cache_tag__T_56_mask) begin
      cache_tag[cache_tag__T_56_addr] <= cache_tag__T_56_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_57_en & cache_tag__T_57_mask) begin
      cache_tag[cache_tag__T_57_addr] <= cache_tag__T_57_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_58_en & cache_tag__T_58_mask) begin
      cache_tag[cache_tag__T_58_addr] <= cache_tag__T_58_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_59_en & cache_tag__T_59_mask) begin
      cache_tag[cache_tag__T_59_addr] <= cache_tag__T_59_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_60_en & cache_tag__T_60_mask) begin
      cache_tag[cache_tag__T_60_addr] <= cache_tag__T_60_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_61_en & cache_tag__T_61_mask) begin
      cache_tag[cache_tag__T_61_addr] <= cache_tag__T_61_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_62_en & cache_tag__T_62_mask) begin
      cache_tag[cache_tag__T_62_addr] <= cache_tag__T_62_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_63_en & cache_tag__T_63_mask) begin
      cache_tag[cache_tag__T_63_addr] <= cache_tag__T_63_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_64_en & cache_tag__T_64_mask) begin
      cache_tag[cache_tag__T_64_addr] <= cache_tag__T_64_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_65_en & cache_tag__T_65_mask) begin
      cache_tag[cache_tag__T_65_addr] <= cache_tag__T_65_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_66_en & cache_tag__T_66_mask) begin
      cache_tag[cache_tag__T_66_addr] <= cache_tag__T_66_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_67_en & cache_tag__T_67_mask) begin
      cache_tag[cache_tag__T_67_addr] <= cache_tag__T_67_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_68_en & cache_tag__T_68_mask) begin
      cache_tag[cache_tag__T_68_addr] <= cache_tag__T_68_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_69_en & cache_tag__T_69_mask) begin
      cache_tag[cache_tag__T_69_addr] <= cache_tag__T_69_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_70_en & cache_tag__T_70_mask) begin
      cache_tag[cache_tag__T_70_addr] <= cache_tag__T_70_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_71_en & cache_tag__T_71_mask) begin
      cache_tag[cache_tag__T_71_addr] <= cache_tag__T_71_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_72_en & cache_tag__T_72_mask) begin
      cache_tag[cache_tag__T_72_addr] <= cache_tag__T_72_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_73_en & cache_tag__T_73_mask) begin
      cache_tag[cache_tag__T_73_addr] <= cache_tag__T_73_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_74_en & cache_tag__T_74_mask) begin
      cache_tag[cache_tag__T_74_addr] <= cache_tag__T_74_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_75_en & cache_tag__T_75_mask) begin
      cache_tag[cache_tag__T_75_addr] <= cache_tag__T_75_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_76_en & cache_tag__T_76_mask) begin
      cache_tag[cache_tag__T_76_addr] <= cache_tag__T_76_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_77_en & cache_tag__T_77_mask) begin
      cache_tag[cache_tag__T_77_addr] <= cache_tag__T_77_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_78_en & cache_tag__T_78_mask) begin
      cache_tag[cache_tag__T_78_addr] <= cache_tag__T_78_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_79_en & cache_tag__T_79_mask) begin
      cache_tag[cache_tag__T_79_addr] <= cache_tag__T_79_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_80_en & cache_tag__T_80_mask) begin
      cache_tag[cache_tag__T_80_addr] <= cache_tag__T_80_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_81_en & cache_tag__T_81_mask) begin
      cache_tag[cache_tag__T_81_addr] <= cache_tag__T_81_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_82_en & cache_tag__T_82_mask) begin
      cache_tag[cache_tag__T_82_addr] <= cache_tag__T_82_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_83_en & cache_tag__T_83_mask) begin
      cache_tag[cache_tag__T_83_addr] <= cache_tag__T_83_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_84_en & cache_tag__T_84_mask) begin
      cache_tag[cache_tag__T_84_addr] <= cache_tag__T_84_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_85_en & cache_tag__T_85_mask) begin
      cache_tag[cache_tag__T_85_addr] <= cache_tag__T_85_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_86_en & cache_tag__T_86_mask) begin
      cache_tag[cache_tag__T_86_addr] <= cache_tag__T_86_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_87_en & cache_tag__T_87_mask) begin
      cache_tag[cache_tag__T_87_addr] <= cache_tag__T_87_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_88_en & cache_tag__T_88_mask) begin
      cache_tag[cache_tag__T_88_addr] <= cache_tag__T_88_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_89_en & cache_tag__T_89_mask) begin
      cache_tag[cache_tag__T_89_addr] <= cache_tag__T_89_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_90_en & cache_tag__T_90_mask) begin
      cache_tag[cache_tag__T_90_addr] <= cache_tag__T_90_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_91_en & cache_tag__T_91_mask) begin
      cache_tag[cache_tag__T_91_addr] <= cache_tag__T_91_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_92_en & cache_tag__T_92_mask) begin
      cache_tag[cache_tag__T_92_addr] <= cache_tag__T_92_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_93_en & cache_tag__T_93_mask) begin
      cache_tag[cache_tag__T_93_addr] <= cache_tag__T_93_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_94_en & cache_tag__T_94_mask) begin
      cache_tag[cache_tag__T_94_addr] <= cache_tag__T_94_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_95_en & cache_tag__T_95_mask) begin
      cache_tag[cache_tag__T_95_addr] <= cache_tag__T_95_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_96_en & cache_tag__T_96_mask) begin
      cache_tag[cache_tag__T_96_addr] <= cache_tag__T_96_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_97_en & cache_tag__T_97_mask) begin
      cache_tag[cache_tag__T_97_addr] <= cache_tag__T_97_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_98_en & cache_tag__T_98_mask) begin
      cache_tag[cache_tag__T_98_addr] <= cache_tag__T_98_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_99_en & cache_tag__T_99_mask) begin
      cache_tag[cache_tag__T_99_addr] <= cache_tag__T_99_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_100_en & cache_tag__T_100_mask) begin
      cache_tag[cache_tag__T_100_addr] <= cache_tag__T_100_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_101_en & cache_tag__T_101_mask) begin
      cache_tag[cache_tag__T_101_addr] <= cache_tag__T_101_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_102_en & cache_tag__T_102_mask) begin
      cache_tag[cache_tag__T_102_addr] <= cache_tag__T_102_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_103_en & cache_tag__T_103_mask) begin
      cache_tag[cache_tag__T_103_addr] <= cache_tag__T_103_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_104_en & cache_tag__T_104_mask) begin
      cache_tag[cache_tag__T_104_addr] <= cache_tag__T_104_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_105_en & cache_tag__T_105_mask) begin
      cache_tag[cache_tag__T_105_addr] <= cache_tag__T_105_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_106_en & cache_tag__T_106_mask) begin
      cache_tag[cache_tag__T_106_addr] <= cache_tag__T_106_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_107_en & cache_tag__T_107_mask) begin
      cache_tag[cache_tag__T_107_addr] <= cache_tag__T_107_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_108_en & cache_tag__T_108_mask) begin
      cache_tag[cache_tag__T_108_addr] <= cache_tag__T_108_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_109_en & cache_tag__T_109_mask) begin
      cache_tag[cache_tag__T_109_addr] <= cache_tag__T_109_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_110_en & cache_tag__T_110_mask) begin
      cache_tag[cache_tag__T_110_addr] <= cache_tag__T_110_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_111_en & cache_tag__T_111_mask) begin
      cache_tag[cache_tag__T_111_addr] <= cache_tag__T_111_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_112_en & cache_tag__T_112_mask) begin
      cache_tag[cache_tag__T_112_addr] <= cache_tag__T_112_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_113_en & cache_tag__T_113_mask) begin
      cache_tag[cache_tag__T_113_addr] <= cache_tag__T_113_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_114_en & cache_tag__T_114_mask) begin
      cache_tag[cache_tag__T_114_addr] <= cache_tag__T_114_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_115_en & cache_tag__T_115_mask) begin
      cache_tag[cache_tag__T_115_addr] <= cache_tag__T_115_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_116_en & cache_tag__T_116_mask) begin
      cache_tag[cache_tag__T_116_addr] <= cache_tag__T_116_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_117_en & cache_tag__T_117_mask) begin
      cache_tag[cache_tag__T_117_addr] <= cache_tag__T_117_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_118_en & cache_tag__T_118_mask) begin
      cache_tag[cache_tag__T_118_addr] <= cache_tag__T_118_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_119_en & cache_tag__T_119_mask) begin
      cache_tag[cache_tag__T_119_addr] <= cache_tag__T_119_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_120_en & cache_tag__T_120_mask) begin
      cache_tag[cache_tag__T_120_addr] <= cache_tag__T_120_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_121_en & cache_tag__T_121_mask) begin
      cache_tag[cache_tag__T_121_addr] <= cache_tag__T_121_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_122_en & cache_tag__T_122_mask) begin
      cache_tag[cache_tag__T_122_addr] <= cache_tag__T_122_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_123_en & cache_tag__T_123_mask) begin
      cache_tag[cache_tag__T_123_addr] <= cache_tag__T_123_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_124_en & cache_tag__T_124_mask) begin
      cache_tag[cache_tag__T_124_addr] <= cache_tag__T_124_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_125_en & cache_tag__T_125_mask) begin
      cache_tag[cache_tag__T_125_addr] <= cache_tag__T_125_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_126_en & cache_tag__T_126_mask) begin
      cache_tag[cache_tag__T_126_addr] <= cache_tag__T_126_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_127_en & cache_tag__T_127_mask) begin
      cache_tag[cache_tag__T_127_addr] <= cache_tag__T_127_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_128_en & cache_tag__T_128_mask) begin
      cache_tag[cache_tag__T_128_addr] <= cache_tag__T_128_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_129_en & cache_tag__T_129_mask) begin
      cache_tag[cache_tag__T_129_addr] <= cache_tag__T_129_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_130_en & cache_tag__T_130_mask) begin
      cache_tag[cache_tag__T_130_addr] <= cache_tag__T_130_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_131_en & cache_tag__T_131_mask) begin
      cache_tag[cache_tag__T_131_addr] <= cache_tag__T_131_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_132_en & cache_tag__T_132_mask) begin
      cache_tag[cache_tag__T_132_addr] <= cache_tag__T_132_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_133_en & cache_tag__T_133_mask) begin
      cache_tag[cache_tag__T_133_addr] <= cache_tag__T_133_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_134_en & cache_tag__T_134_mask) begin
      cache_tag[cache_tag__T_134_addr] <= cache_tag__T_134_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_135_en & cache_tag__T_135_mask) begin
      cache_tag[cache_tag__T_135_addr] <= cache_tag__T_135_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_136_en & cache_tag__T_136_mask) begin
      cache_tag[cache_tag__T_136_addr] <= cache_tag__T_136_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_137_en & cache_tag__T_137_mask) begin
      cache_tag[cache_tag__T_137_addr] <= cache_tag__T_137_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_138_en & cache_tag__T_138_mask) begin
      cache_tag[cache_tag__T_138_addr] <= cache_tag__T_138_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_139_en & cache_tag__T_139_mask) begin
      cache_tag[cache_tag__T_139_addr] <= cache_tag__T_139_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_140_en & cache_tag__T_140_mask) begin
      cache_tag[cache_tag__T_140_addr] <= cache_tag__T_140_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_141_en & cache_tag__T_141_mask) begin
      cache_tag[cache_tag__T_141_addr] <= cache_tag__T_141_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_142_en & cache_tag__T_142_mask) begin
      cache_tag[cache_tag__T_142_addr] <= cache_tag__T_142_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_143_en & cache_tag__T_143_mask) begin
      cache_tag[cache_tag__T_143_addr] <= cache_tag__T_143_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_144_en & cache_tag__T_144_mask) begin
      cache_tag[cache_tag__T_144_addr] <= cache_tag__T_144_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_145_en & cache_tag__T_145_mask) begin
      cache_tag[cache_tag__T_145_addr] <= cache_tag__T_145_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_146_en & cache_tag__T_146_mask) begin
      cache_tag[cache_tag__T_146_addr] <= cache_tag__T_146_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_147_en & cache_tag__T_147_mask) begin
      cache_tag[cache_tag__T_147_addr] <= cache_tag__T_147_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_148_en & cache_tag__T_148_mask) begin
      cache_tag[cache_tag__T_148_addr] <= cache_tag__T_148_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_149_en & cache_tag__T_149_mask) begin
      cache_tag[cache_tag__T_149_addr] <= cache_tag__T_149_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_150_en & cache_tag__T_150_mask) begin
      cache_tag[cache_tag__T_150_addr] <= cache_tag__T_150_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_151_en & cache_tag__T_151_mask) begin
      cache_tag[cache_tag__T_151_addr] <= cache_tag__T_151_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_152_en & cache_tag__T_152_mask) begin
      cache_tag[cache_tag__T_152_addr] <= cache_tag__T_152_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_153_en & cache_tag__T_153_mask) begin
      cache_tag[cache_tag__T_153_addr] <= cache_tag__T_153_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_154_en & cache_tag__T_154_mask) begin
      cache_tag[cache_tag__T_154_addr] <= cache_tag__T_154_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_155_en & cache_tag__T_155_mask) begin
      cache_tag[cache_tag__T_155_addr] <= cache_tag__T_155_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_156_en & cache_tag__T_156_mask) begin
      cache_tag[cache_tag__T_156_addr] <= cache_tag__T_156_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_157_en & cache_tag__T_157_mask) begin
      cache_tag[cache_tag__T_157_addr] <= cache_tag__T_157_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_158_en & cache_tag__T_158_mask) begin
      cache_tag[cache_tag__T_158_addr] <= cache_tag__T_158_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_159_en & cache_tag__T_159_mask) begin
      cache_tag[cache_tag__T_159_addr] <= cache_tag__T_159_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_160_en & cache_tag__T_160_mask) begin
      cache_tag[cache_tag__T_160_addr] <= cache_tag__T_160_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_161_en & cache_tag__T_161_mask) begin
      cache_tag[cache_tag__T_161_addr] <= cache_tag__T_161_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_162_en & cache_tag__T_162_mask) begin
      cache_tag[cache_tag__T_162_addr] <= cache_tag__T_162_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_163_en & cache_tag__T_163_mask) begin
      cache_tag[cache_tag__T_163_addr] <= cache_tag__T_163_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_164_en & cache_tag__T_164_mask) begin
      cache_tag[cache_tag__T_164_addr] <= cache_tag__T_164_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_165_en & cache_tag__T_165_mask) begin
      cache_tag[cache_tag__T_165_addr] <= cache_tag__T_165_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_166_en & cache_tag__T_166_mask) begin
      cache_tag[cache_tag__T_166_addr] <= cache_tag__T_166_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_167_en & cache_tag__T_167_mask) begin
      cache_tag[cache_tag__T_167_addr] <= cache_tag__T_167_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_168_en & cache_tag__T_168_mask) begin
      cache_tag[cache_tag__T_168_addr] <= cache_tag__T_168_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_169_en & cache_tag__T_169_mask) begin
      cache_tag[cache_tag__T_169_addr] <= cache_tag__T_169_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_170_en & cache_tag__T_170_mask) begin
      cache_tag[cache_tag__T_170_addr] <= cache_tag__T_170_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_171_en & cache_tag__T_171_mask) begin
      cache_tag[cache_tag__T_171_addr] <= cache_tag__T_171_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_172_en & cache_tag__T_172_mask) begin
      cache_tag[cache_tag__T_172_addr] <= cache_tag__T_172_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_173_en & cache_tag__T_173_mask) begin
      cache_tag[cache_tag__T_173_addr] <= cache_tag__T_173_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_174_en & cache_tag__T_174_mask) begin
      cache_tag[cache_tag__T_174_addr] <= cache_tag__T_174_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_175_en & cache_tag__T_175_mask) begin
      cache_tag[cache_tag__T_175_addr] <= cache_tag__T_175_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_176_en & cache_tag__T_176_mask) begin
      cache_tag[cache_tag__T_176_addr] <= cache_tag__T_176_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_177_en & cache_tag__T_177_mask) begin
      cache_tag[cache_tag__T_177_addr] <= cache_tag__T_177_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_178_en & cache_tag__T_178_mask) begin
      cache_tag[cache_tag__T_178_addr] <= cache_tag__T_178_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_179_en & cache_tag__T_179_mask) begin
      cache_tag[cache_tag__T_179_addr] <= cache_tag__T_179_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_180_en & cache_tag__T_180_mask) begin
      cache_tag[cache_tag__T_180_addr] <= cache_tag__T_180_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_181_en & cache_tag__T_181_mask) begin
      cache_tag[cache_tag__T_181_addr] <= cache_tag__T_181_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_182_en & cache_tag__T_182_mask) begin
      cache_tag[cache_tag__T_182_addr] <= cache_tag__T_182_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_183_en & cache_tag__T_183_mask) begin
      cache_tag[cache_tag__T_183_addr] <= cache_tag__T_183_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_184_en & cache_tag__T_184_mask) begin
      cache_tag[cache_tag__T_184_addr] <= cache_tag__T_184_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_185_en & cache_tag__T_185_mask) begin
      cache_tag[cache_tag__T_185_addr] <= cache_tag__T_185_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_186_en & cache_tag__T_186_mask) begin
      cache_tag[cache_tag__T_186_addr] <= cache_tag__T_186_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_187_en & cache_tag__T_187_mask) begin
      cache_tag[cache_tag__T_187_addr] <= cache_tag__T_187_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_188_en & cache_tag__T_188_mask) begin
      cache_tag[cache_tag__T_188_addr] <= cache_tag__T_188_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_189_en & cache_tag__T_189_mask) begin
      cache_tag[cache_tag__T_189_addr] <= cache_tag__T_189_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_190_en & cache_tag__T_190_mask) begin
      cache_tag[cache_tag__T_190_addr] <= cache_tag__T_190_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_191_en & cache_tag__T_191_mask) begin
      cache_tag[cache_tag__T_191_addr] <= cache_tag__T_191_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_192_en & cache_tag__T_192_mask) begin
      cache_tag[cache_tag__T_192_addr] <= cache_tag__T_192_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_193_en & cache_tag__T_193_mask) begin
      cache_tag[cache_tag__T_193_addr] <= cache_tag__T_193_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_194_en & cache_tag__T_194_mask) begin
      cache_tag[cache_tag__T_194_addr] <= cache_tag__T_194_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_195_en & cache_tag__T_195_mask) begin
      cache_tag[cache_tag__T_195_addr] <= cache_tag__T_195_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_196_en & cache_tag__T_196_mask) begin
      cache_tag[cache_tag__T_196_addr] <= cache_tag__T_196_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_197_en & cache_tag__T_197_mask) begin
      cache_tag[cache_tag__T_197_addr] <= cache_tag__T_197_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_198_en & cache_tag__T_198_mask) begin
      cache_tag[cache_tag__T_198_addr] <= cache_tag__T_198_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_199_en & cache_tag__T_199_mask) begin
      cache_tag[cache_tag__T_199_addr] <= cache_tag__T_199_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_200_en & cache_tag__T_200_mask) begin
      cache_tag[cache_tag__T_200_addr] <= cache_tag__T_200_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_201_en & cache_tag__T_201_mask) begin
      cache_tag[cache_tag__T_201_addr] <= cache_tag__T_201_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_202_en & cache_tag__T_202_mask) begin
      cache_tag[cache_tag__T_202_addr] <= cache_tag__T_202_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_203_en & cache_tag__T_203_mask) begin
      cache_tag[cache_tag__T_203_addr] <= cache_tag__T_203_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_204_en & cache_tag__T_204_mask) begin
      cache_tag[cache_tag__T_204_addr] <= cache_tag__T_204_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_205_en & cache_tag__T_205_mask) begin
      cache_tag[cache_tag__T_205_addr] <= cache_tag__T_205_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_206_en & cache_tag__T_206_mask) begin
      cache_tag[cache_tag__T_206_addr] <= cache_tag__T_206_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_207_en & cache_tag__T_207_mask) begin
      cache_tag[cache_tag__T_207_addr] <= cache_tag__T_207_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_208_en & cache_tag__T_208_mask) begin
      cache_tag[cache_tag__T_208_addr] <= cache_tag__T_208_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_209_en & cache_tag__T_209_mask) begin
      cache_tag[cache_tag__T_209_addr] <= cache_tag__T_209_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_210_en & cache_tag__T_210_mask) begin
      cache_tag[cache_tag__T_210_addr] <= cache_tag__T_210_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_211_en & cache_tag__T_211_mask) begin
      cache_tag[cache_tag__T_211_addr] <= cache_tag__T_211_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_212_en & cache_tag__T_212_mask) begin
      cache_tag[cache_tag__T_212_addr] <= cache_tag__T_212_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_213_en & cache_tag__T_213_mask) begin
      cache_tag[cache_tag__T_213_addr] <= cache_tag__T_213_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_214_en & cache_tag__T_214_mask) begin
      cache_tag[cache_tag__T_214_addr] <= cache_tag__T_214_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_215_en & cache_tag__T_215_mask) begin
      cache_tag[cache_tag__T_215_addr] <= cache_tag__T_215_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_216_en & cache_tag__T_216_mask) begin
      cache_tag[cache_tag__T_216_addr] <= cache_tag__T_216_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_217_en & cache_tag__T_217_mask) begin
      cache_tag[cache_tag__T_217_addr] <= cache_tag__T_217_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_218_en & cache_tag__T_218_mask) begin
      cache_tag[cache_tag__T_218_addr] <= cache_tag__T_218_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_219_en & cache_tag__T_219_mask) begin
      cache_tag[cache_tag__T_219_addr] <= cache_tag__T_219_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_220_en & cache_tag__T_220_mask) begin
      cache_tag[cache_tag__T_220_addr] <= cache_tag__T_220_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_221_en & cache_tag__T_221_mask) begin
      cache_tag[cache_tag__T_221_addr] <= cache_tag__T_221_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_222_en & cache_tag__T_222_mask) begin
      cache_tag[cache_tag__T_222_addr] <= cache_tag__T_222_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_223_en & cache_tag__T_223_mask) begin
      cache_tag[cache_tag__T_223_addr] <= cache_tag__T_223_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_224_en & cache_tag__T_224_mask) begin
      cache_tag[cache_tag__T_224_addr] <= cache_tag__T_224_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_225_en & cache_tag__T_225_mask) begin
      cache_tag[cache_tag__T_225_addr] <= cache_tag__T_225_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_226_en & cache_tag__T_226_mask) begin
      cache_tag[cache_tag__T_226_addr] <= cache_tag__T_226_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_227_en & cache_tag__T_227_mask) begin
      cache_tag[cache_tag__T_227_addr] <= cache_tag__T_227_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_228_en & cache_tag__T_228_mask) begin
      cache_tag[cache_tag__T_228_addr] <= cache_tag__T_228_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_229_en & cache_tag__T_229_mask) begin
      cache_tag[cache_tag__T_229_addr] <= cache_tag__T_229_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_230_en & cache_tag__T_230_mask) begin
      cache_tag[cache_tag__T_230_addr] <= cache_tag__T_230_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_231_en & cache_tag__T_231_mask) begin
      cache_tag[cache_tag__T_231_addr] <= cache_tag__T_231_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_232_en & cache_tag__T_232_mask) begin
      cache_tag[cache_tag__T_232_addr] <= cache_tag__T_232_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_233_en & cache_tag__T_233_mask) begin
      cache_tag[cache_tag__T_233_addr] <= cache_tag__T_233_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_234_en & cache_tag__T_234_mask) begin
      cache_tag[cache_tag__T_234_addr] <= cache_tag__T_234_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_235_en & cache_tag__T_235_mask) begin
      cache_tag[cache_tag__T_235_addr] <= cache_tag__T_235_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_236_en & cache_tag__T_236_mask) begin
      cache_tag[cache_tag__T_236_addr] <= cache_tag__T_236_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_237_en & cache_tag__T_237_mask) begin
      cache_tag[cache_tag__T_237_addr] <= cache_tag__T_237_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_238_en & cache_tag__T_238_mask) begin
      cache_tag[cache_tag__T_238_addr] <= cache_tag__T_238_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_239_en & cache_tag__T_239_mask) begin
      cache_tag[cache_tag__T_239_addr] <= cache_tag__T_239_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_240_en & cache_tag__T_240_mask) begin
      cache_tag[cache_tag__T_240_addr] <= cache_tag__T_240_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_241_en & cache_tag__T_241_mask) begin
      cache_tag[cache_tag__T_241_addr] <= cache_tag__T_241_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_242_en & cache_tag__T_242_mask) begin
      cache_tag[cache_tag__T_242_addr] <= cache_tag__T_242_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_243_en & cache_tag__T_243_mask) begin
      cache_tag[cache_tag__T_243_addr] <= cache_tag__T_243_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_244_en & cache_tag__T_244_mask) begin
      cache_tag[cache_tag__T_244_addr] <= cache_tag__T_244_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_245_en & cache_tag__T_245_mask) begin
      cache_tag[cache_tag__T_245_addr] <= cache_tag__T_245_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_246_en & cache_tag__T_246_mask) begin
      cache_tag[cache_tag__T_246_addr] <= cache_tag__T_246_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_247_en & cache_tag__T_247_mask) begin
      cache_tag[cache_tag__T_247_addr] <= cache_tag__T_247_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_248_en & cache_tag__T_248_mask) begin
      cache_tag[cache_tag__T_248_addr] <= cache_tag__T_248_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_249_en & cache_tag__T_249_mask) begin
      cache_tag[cache_tag__T_249_addr] <= cache_tag__T_249_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_250_en & cache_tag__T_250_mask) begin
      cache_tag[cache_tag__T_250_addr] <= cache_tag__T_250_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_251_en & cache_tag__T_251_mask) begin
      cache_tag[cache_tag__T_251_addr] <= cache_tag__T_251_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_252_en & cache_tag__T_252_mask) begin
      cache_tag[cache_tag__T_252_addr] <= cache_tag__T_252_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_253_en & cache_tag__T_253_mask) begin
      cache_tag[cache_tag__T_253_addr] <= cache_tag__T_253_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_254_en & cache_tag__T_254_mask) begin
      cache_tag[cache_tag__T_254_addr] <= cache_tag__T_254_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_255_en & cache_tag__T_255_mask) begin
      cache_tag[cache_tag__T_255_addr] <= cache_tag__T_255_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_256_en & cache_tag__T_256_mask) begin
      cache_tag[cache_tag__T_256_addr] <= cache_tag__T_256_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_257_en & cache_tag__T_257_mask) begin
      cache_tag[cache_tag__T_257_addr] <= cache_tag__T_257_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_258_en & cache_tag__T_258_mask) begin
      cache_tag[cache_tag__T_258_addr] <= cache_tag__T_258_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_259_en & cache_tag__T_259_mask) begin
      cache_tag[cache_tag__T_259_addr] <= cache_tag__T_259_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_260_en & cache_tag__T_260_mask) begin
      cache_tag[cache_tag__T_260_addr] <= cache_tag__T_260_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_261_en & cache_tag__T_261_mask) begin
      cache_tag[cache_tag__T_261_addr] <= cache_tag__T_261_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_262_en & cache_tag__T_262_mask) begin
      cache_tag[cache_tag__T_262_addr] <= cache_tag__T_262_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_263_en & cache_tag__T_263_mask) begin
      cache_tag[cache_tag__T_263_addr] <= cache_tag__T_263_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_264_en & cache_tag__T_264_mask) begin
      cache_tag[cache_tag__T_264_addr] <= cache_tag__T_264_data; // @[icache.scala 91:18]
    end
    if(cache_tag__T_265_en & cache_tag__T_265_mask) begin
      cache_tag[cache_tag__T_265_addr] <= cache_tag__T_265_data; // @[icache.scala 91:18]
    end
    if(cache_tag_s1_entry_w_en & cache_tag_s1_entry_w_mask) begin
      cache_tag[cache_tag_s1_entry_w_addr] <= cache_tag_s1_entry_w_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_8_en & cache_data__T_8_mask) begin
      cache_data[cache_data__T_8_addr] <= cache_data__T_8_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_10_en & cache_data__T_10_mask) begin
      cache_data[cache_data__T_10_addr] <= cache_data__T_10_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_11_en & cache_data__T_11_mask) begin
      cache_data[cache_data__T_11_addr] <= cache_data__T_11_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_12_en & cache_data__T_12_mask) begin
      cache_data[cache_data__T_12_addr] <= cache_data__T_12_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_13_en & cache_data__T_13_mask) begin
      cache_data[cache_data__T_13_addr] <= cache_data__T_13_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_14_en & cache_data__T_14_mask) begin
      cache_data[cache_data__T_14_addr] <= cache_data__T_14_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_15_en & cache_data__T_15_mask) begin
      cache_data[cache_data__T_15_addr] <= cache_data__T_15_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_16_en & cache_data__T_16_mask) begin
      cache_data[cache_data__T_16_addr] <= cache_data__T_16_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_17_en & cache_data__T_17_mask) begin
      cache_data[cache_data__T_17_addr] <= cache_data__T_17_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_18_en & cache_data__T_18_mask) begin
      cache_data[cache_data__T_18_addr] <= cache_data__T_18_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_19_en & cache_data__T_19_mask) begin
      cache_data[cache_data__T_19_addr] <= cache_data__T_19_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_20_en & cache_data__T_20_mask) begin
      cache_data[cache_data__T_20_addr] <= cache_data__T_20_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_21_en & cache_data__T_21_mask) begin
      cache_data[cache_data__T_21_addr] <= cache_data__T_21_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_22_en & cache_data__T_22_mask) begin
      cache_data[cache_data__T_22_addr] <= cache_data__T_22_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_23_en & cache_data__T_23_mask) begin
      cache_data[cache_data__T_23_addr] <= cache_data__T_23_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_24_en & cache_data__T_24_mask) begin
      cache_data[cache_data__T_24_addr] <= cache_data__T_24_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_25_en & cache_data__T_25_mask) begin
      cache_data[cache_data__T_25_addr] <= cache_data__T_25_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_26_en & cache_data__T_26_mask) begin
      cache_data[cache_data__T_26_addr] <= cache_data__T_26_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_27_en & cache_data__T_27_mask) begin
      cache_data[cache_data__T_27_addr] <= cache_data__T_27_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_28_en & cache_data__T_28_mask) begin
      cache_data[cache_data__T_28_addr] <= cache_data__T_28_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_29_en & cache_data__T_29_mask) begin
      cache_data[cache_data__T_29_addr] <= cache_data__T_29_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_30_en & cache_data__T_30_mask) begin
      cache_data[cache_data__T_30_addr] <= cache_data__T_30_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_31_en & cache_data__T_31_mask) begin
      cache_data[cache_data__T_31_addr] <= cache_data__T_31_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_32_en & cache_data__T_32_mask) begin
      cache_data[cache_data__T_32_addr] <= cache_data__T_32_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_33_en & cache_data__T_33_mask) begin
      cache_data[cache_data__T_33_addr] <= cache_data__T_33_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_34_en & cache_data__T_34_mask) begin
      cache_data[cache_data__T_34_addr] <= cache_data__T_34_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_35_en & cache_data__T_35_mask) begin
      cache_data[cache_data__T_35_addr] <= cache_data__T_35_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_36_en & cache_data__T_36_mask) begin
      cache_data[cache_data__T_36_addr] <= cache_data__T_36_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_37_en & cache_data__T_37_mask) begin
      cache_data[cache_data__T_37_addr] <= cache_data__T_37_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_38_en & cache_data__T_38_mask) begin
      cache_data[cache_data__T_38_addr] <= cache_data__T_38_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_39_en & cache_data__T_39_mask) begin
      cache_data[cache_data__T_39_addr] <= cache_data__T_39_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_40_en & cache_data__T_40_mask) begin
      cache_data[cache_data__T_40_addr] <= cache_data__T_40_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_41_en & cache_data__T_41_mask) begin
      cache_data[cache_data__T_41_addr] <= cache_data__T_41_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_42_en & cache_data__T_42_mask) begin
      cache_data[cache_data__T_42_addr] <= cache_data__T_42_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_43_en & cache_data__T_43_mask) begin
      cache_data[cache_data__T_43_addr] <= cache_data__T_43_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_44_en & cache_data__T_44_mask) begin
      cache_data[cache_data__T_44_addr] <= cache_data__T_44_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_45_en & cache_data__T_45_mask) begin
      cache_data[cache_data__T_45_addr] <= cache_data__T_45_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_46_en & cache_data__T_46_mask) begin
      cache_data[cache_data__T_46_addr] <= cache_data__T_46_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_47_en & cache_data__T_47_mask) begin
      cache_data[cache_data__T_47_addr] <= cache_data__T_47_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_48_en & cache_data__T_48_mask) begin
      cache_data[cache_data__T_48_addr] <= cache_data__T_48_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_49_en & cache_data__T_49_mask) begin
      cache_data[cache_data__T_49_addr] <= cache_data__T_49_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_50_en & cache_data__T_50_mask) begin
      cache_data[cache_data__T_50_addr] <= cache_data__T_50_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_51_en & cache_data__T_51_mask) begin
      cache_data[cache_data__T_51_addr] <= cache_data__T_51_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_52_en & cache_data__T_52_mask) begin
      cache_data[cache_data__T_52_addr] <= cache_data__T_52_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_53_en & cache_data__T_53_mask) begin
      cache_data[cache_data__T_53_addr] <= cache_data__T_53_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_54_en & cache_data__T_54_mask) begin
      cache_data[cache_data__T_54_addr] <= cache_data__T_54_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_55_en & cache_data__T_55_mask) begin
      cache_data[cache_data__T_55_addr] <= cache_data__T_55_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_56_en & cache_data__T_56_mask) begin
      cache_data[cache_data__T_56_addr] <= cache_data__T_56_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_57_en & cache_data__T_57_mask) begin
      cache_data[cache_data__T_57_addr] <= cache_data__T_57_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_58_en & cache_data__T_58_mask) begin
      cache_data[cache_data__T_58_addr] <= cache_data__T_58_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_59_en & cache_data__T_59_mask) begin
      cache_data[cache_data__T_59_addr] <= cache_data__T_59_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_60_en & cache_data__T_60_mask) begin
      cache_data[cache_data__T_60_addr] <= cache_data__T_60_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_61_en & cache_data__T_61_mask) begin
      cache_data[cache_data__T_61_addr] <= cache_data__T_61_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_62_en & cache_data__T_62_mask) begin
      cache_data[cache_data__T_62_addr] <= cache_data__T_62_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_63_en & cache_data__T_63_mask) begin
      cache_data[cache_data__T_63_addr] <= cache_data__T_63_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_64_en & cache_data__T_64_mask) begin
      cache_data[cache_data__T_64_addr] <= cache_data__T_64_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_65_en & cache_data__T_65_mask) begin
      cache_data[cache_data__T_65_addr] <= cache_data__T_65_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_66_en & cache_data__T_66_mask) begin
      cache_data[cache_data__T_66_addr] <= cache_data__T_66_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_67_en & cache_data__T_67_mask) begin
      cache_data[cache_data__T_67_addr] <= cache_data__T_67_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_68_en & cache_data__T_68_mask) begin
      cache_data[cache_data__T_68_addr] <= cache_data__T_68_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_69_en & cache_data__T_69_mask) begin
      cache_data[cache_data__T_69_addr] <= cache_data__T_69_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_70_en & cache_data__T_70_mask) begin
      cache_data[cache_data__T_70_addr] <= cache_data__T_70_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_71_en & cache_data__T_71_mask) begin
      cache_data[cache_data__T_71_addr] <= cache_data__T_71_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_72_en & cache_data__T_72_mask) begin
      cache_data[cache_data__T_72_addr] <= cache_data__T_72_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_73_en & cache_data__T_73_mask) begin
      cache_data[cache_data__T_73_addr] <= cache_data__T_73_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_74_en & cache_data__T_74_mask) begin
      cache_data[cache_data__T_74_addr] <= cache_data__T_74_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_75_en & cache_data__T_75_mask) begin
      cache_data[cache_data__T_75_addr] <= cache_data__T_75_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_76_en & cache_data__T_76_mask) begin
      cache_data[cache_data__T_76_addr] <= cache_data__T_76_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_77_en & cache_data__T_77_mask) begin
      cache_data[cache_data__T_77_addr] <= cache_data__T_77_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_78_en & cache_data__T_78_mask) begin
      cache_data[cache_data__T_78_addr] <= cache_data__T_78_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_79_en & cache_data__T_79_mask) begin
      cache_data[cache_data__T_79_addr] <= cache_data__T_79_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_80_en & cache_data__T_80_mask) begin
      cache_data[cache_data__T_80_addr] <= cache_data__T_80_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_81_en & cache_data__T_81_mask) begin
      cache_data[cache_data__T_81_addr] <= cache_data__T_81_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_82_en & cache_data__T_82_mask) begin
      cache_data[cache_data__T_82_addr] <= cache_data__T_82_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_83_en & cache_data__T_83_mask) begin
      cache_data[cache_data__T_83_addr] <= cache_data__T_83_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_84_en & cache_data__T_84_mask) begin
      cache_data[cache_data__T_84_addr] <= cache_data__T_84_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_85_en & cache_data__T_85_mask) begin
      cache_data[cache_data__T_85_addr] <= cache_data__T_85_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_86_en & cache_data__T_86_mask) begin
      cache_data[cache_data__T_86_addr] <= cache_data__T_86_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_87_en & cache_data__T_87_mask) begin
      cache_data[cache_data__T_87_addr] <= cache_data__T_87_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_88_en & cache_data__T_88_mask) begin
      cache_data[cache_data__T_88_addr] <= cache_data__T_88_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_89_en & cache_data__T_89_mask) begin
      cache_data[cache_data__T_89_addr] <= cache_data__T_89_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_90_en & cache_data__T_90_mask) begin
      cache_data[cache_data__T_90_addr] <= cache_data__T_90_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_91_en & cache_data__T_91_mask) begin
      cache_data[cache_data__T_91_addr] <= cache_data__T_91_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_92_en & cache_data__T_92_mask) begin
      cache_data[cache_data__T_92_addr] <= cache_data__T_92_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_93_en & cache_data__T_93_mask) begin
      cache_data[cache_data__T_93_addr] <= cache_data__T_93_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_94_en & cache_data__T_94_mask) begin
      cache_data[cache_data__T_94_addr] <= cache_data__T_94_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_95_en & cache_data__T_95_mask) begin
      cache_data[cache_data__T_95_addr] <= cache_data__T_95_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_96_en & cache_data__T_96_mask) begin
      cache_data[cache_data__T_96_addr] <= cache_data__T_96_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_97_en & cache_data__T_97_mask) begin
      cache_data[cache_data__T_97_addr] <= cache_data__T_97_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_98_en & cache_data__T_98_mask) begin
      cache_data[cache_data__T_98_addr] <= cache_data__T_98_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_99_en & cache_data__T_99_mask) begin
      cache_data[cache_data__T_99_addr] <= cache_data__T_99_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_100_en & cache_data__T_100_mask) begin
      cache_data[cache_data__T_100_addr] <= cache_data__T_100_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_101_en & cache_data__T_101_mask) begin
      cache_data[cache_data__T_101_addr] <= cache_data__T_101_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_102_en & cache_data__T_102_mask) begin
      cache_data[cache_data__T_102_addr] <= cache_data__T_102_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_103_en & cache_data__T_103_mask) begin
      cache_data[cache_data__T_103_addr] <= cache_data__T_103_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_104_en & cache_data__T_104_mask) begin
      cache_data[cache_data__T_104_addr] <= cache_data__T_104_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_105_en & cache_data__T_105_mask) begin
      cache_data[cache_data__T_105_addr] <= cache_data__T_105_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_106_en & cache_data__T_106_mask) begin
      cache_data[cache_data__T_106_addr] <= cache_data__T_106_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_107_en & cache_data__T_107_mask) begin
      cache_data[cache_data__T_107_addr] <= cache_data__T_107_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_108_en & cache_data__T_108_mask) begin
      cache_data[cache_data__T_108_addr] <= cache_data__T_108_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_109_en & cache_data__T_109_mask) begin
      cache_data[cache_data__T_109_addr] <= cache_data__T_109_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_110_en & cache_data__T_110_mask) begin
      cache_data[cache_data__T_110_addr] <= cache_data__T_110_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_111_en & cache_data__T_111_mask) begin
      cache_data[cache_data__T_111_addr] <= cache_data__T_111_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_112_en & cache_data__T_112_mask) begin
      cache_data[cache_data__T_112_addr] <= cache_data__T_112_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_113_en & cache_data__T_113_mask) begin
      cache_data[cache_data__T_113_addr] <= cache_data__T_113_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_114_en & cache_data__T_114_mask) begin
      cache_data[cache_data__T_114_addr] <= cache_data__T_114_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_115_en & cache_data__T_115_mask) begin
      cache_data[cache_data__T_115_addr] <= cache_data__T_115_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_116_en & cache_data__T_116_mask) begin
      cache_data[cache_data__T_116_addr] <= cache_data__T_116_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_117_en & cache_data__T_117_mask) begin
      cache_data[cache_data__T_117_addr] <= cache_data__T_117_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_118_en & cache_data__T_118_mask) begin
      cache_data[cache_data__T_118_addr] <= cache_data__T_118_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_119_en & cache_data__T_119_mask) begin
      cache_data[cache_data__T_119_addr] <= cache_data__T_119_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_120_en & cache_data__T_120_mask) begin
      cache_data[cache_data__T_120_addr] <= cache_data__T_120_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_121_en & cache_data__T_121_mask) begin
      cache_data[cache_data__T_121_addr] <= cache_data__T_121_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_122_en & cache_data__T_122_mask) begin
      cache_data[cache_data__T_122_addr] <= cache_data__T_122_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_123_en & cache_data__T_123_mask) begin
      cache_data[cache_data__T_123_addr] <= cache_data__T_123_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_124_en & cache_data__T_124_mask) begin
      cache_data[cache_data__T_124_addr] <= cache_data__T_124_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_125_en & cache_data__T_125_mask) begin
      cache_data[cache_data__T_125_addr] <= cache_data__T_125_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_126_en & cache_data__T_126_mask) begin
      cache_data[cache_data__T_126_addr] <= cache_data__T_126_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_127_en & cache_data__T_127_mask) begin
      cache_data[cache_data__T_127_addr] <= cache_data__T_127_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_128_en & cache_data__T_128_mask) begin
      cache_data[cache_data__T_128_addr] <= cache_data__T_128_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_129_en & cache_data__T_129_mask) begin
      cache_data[cache_data__T_129_addr] <= cache_data__T_129_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_130_en & cache_data__T_130_mask) begin
      cache_data[cache_data__T_130_addr] <= cache_data__T_130_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_131_en & cache_data__T_131_mask) begin
      cache_data[cache_data__T_131_addr] <= cache_data__T_131_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_132_en & cache_data__T_132_mask) begin
      cache_data[cache_data__T_132_addr] <= cache_data__T_132_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_133_en & cache_data__T_133_mask) begin
      cache_data[cache_data__T_133_addr] <= cache_data__T_133_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_134_en & cache_data__T_134_mask) begin
      cache_data[cache_data__T_134_addr] <= cache_data__T_134_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_135_en & cache_data__T_135_mask) begin
      cache_data[cache_data__T_135_addr] <= cache_data__T_135_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_136_en & cache_data__T_136_mask) begin
      cache_data[cache_data__T_136_addr] <= cache_data__T_136_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_137_en & cache_data__T_137_mask) begin
      cache_data[cache_data__T_137_addr] <= cache_data__T_137_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_138_en & cache_data__T_138_mask) begin
      cache_data[cache_data__T_138_addr] <= cache_data__T_138_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_139_en & cache_data__T_139_mask) begin
      cache_data[cache_data__T_139_addr] <= cache_data__T_139_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_140_en & cache_data__T_140_mask) begin
      cache_data[cache_data__T_140_addr] <= cache_data__T_140_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_141_en & cache_data__T_141_mask) begin
      cache_data[cache_data__T_141_addr] <= cache_data__T_141_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_142_en & cache_data__T_142_mask) begin
      cache_data[cache_data__T_142_addr] <= cache_data__T_142_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_143_en & cache_data__T_143_mask) begin
      cache_data[cache_data__T_143_addr] <= cache_data__T_143_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_144_en & cache_data__T_144_mask) begin
      cache_data[cache_data__T_144_addr] <= cache_data__T_144_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_145_en & cache_data__T_145_mask) begin
      cache_data[cache_data__T_145_addr] <= cache_data__T_145_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_146_en & cache_data__T_146_mask) begin
      cache_data[cache_data__T_146_addr] <= cache_data__T_146_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_147_en & cache_data__T_147_mask) begin
      cache_data[cache_data__T_147_addr] <= cache_data__T_147_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_148_en & cache_data__T_148_mask) begin
      cache_data[cache_data__T_148_addr] <= cache_data__T_148_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_149_en & cache_data__T_149_mask) begin
      cache_data[cache_data__T_149_addr] <= cache_data__T_149_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_150_en & cache_data__T_150_mask) begin
      cache_data[cache_data__T_150_addr] <= cache_data__T_150_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_151_en & cache_data__T_151_mask) begin
      cache_data[cache_data__T_151_addr] <= cache_data__T_151_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_152_en & cache_data__T_152_mask) begin
      cache_data[cache_data__T_152_addr] <= cache_data__T_152_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_153_en & cache_data__T_153_mask) begin
      cache_data[cache_data__T_153_addr] <= cache_data__T_153_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_154_en & cache_data__T_154_mask) begin
      cache_data[cache_data__T_154_addr] <= cache_data__T_154_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_155_en & cache_data__T_155_mask) begin
      cache_data[cache_data__T_155_addr] <= cache_data__T_155_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_156_en & cache_data__T_156_mask) begin
      cache_data[cache_data__T_156_addr] <= cache_data__T_156_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_157_en & cache_data__T_157_mask) begin
      cache_data[cache_data__T_157_addr] <= cache_data__T_157_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_158_en & cache_data__T_158_mask) begin
      cache_data[cache_data__T_158_addr] <= cache_data__T_158_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_159_en & cache_data__T_159_mask) begin
      cache_data[cache_data__T_159_addr] <= cache_data__T_159_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_160_en & cache_data__T_160_mask) begin
      cache_data[cache_data__T_160_addr] <= cache_data__T_160_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_161_en & cache_data__T_161_mask) begin
      cache_data[cache_data__T_161_addr] <= cache_data__T_161_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_162_en & cache_data__T_162_mask) begin
      cache_data[cache_data__T_162_addr] <= cache_data__T_162_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_163_en & cache_data__T_163_mask) begin
      cache_data[cache_data__T_163_addr] <= cache_data__T_163_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_164_en & cache_data__T_164_mask) begin
      cache_data[cache_data__T_164_addr] <= cache_data__T_164_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_165_en & cache_data__T_165_mask) begin
      cache_data[cache_data__T_165_addr] <= cache_data__T_165_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_166_en & cache_data__T_166_mask) begin
      cache_data[cache_data__T_166_addr] <= cache_data__T_166_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_167_en & cache_data__T_167_mask) begin
      cache_data[cache_data__T_167_addr] <= cache_data__T_167_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_168_en & cache_data__T_168_mask) begin
      cache_data[cache_data__T_168_addr] <= cache_data__T_168_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_169_en & cache_data__T_169_mask) begin
      cache_data[cache_data__T_169_addr] <= cache_data__T_169_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_170_en & cache_data__T_170_mask) begin
      cache_data[cache_data__T_170_addr] <= cache_data__T_170_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_171_en & cache_data__T_171_mask) begin
      cache_data[cache_data__T_171_addr] <= cache_data__T_171_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_172_en & cache_data__T_172_mask) begin
      cache_data[cache_data__T_172_addr] <= cache_data__T_172_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_173_en & cache_data__T_173_mask) begin
      cache_data[cache_data__T_173_addr] <= cache_data__T_173_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_174_en & cache_data__T_174_mask) begin
      cache_data[cache_data__T_174_addr] <= cache_data__T_174_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_175_en & cache_data__T_175_mask) begin
      cache_data[cache_data__T_175_addr] <= cache_data__T_175_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_176_en & cache_data__T_176_mask) begin
      cache_data[cache_data__T_176_addr] <= cache_data__T_176_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_177_en & cache_data__T_177_mask) begin
      cache_data[cache_data__T_177_addr] <= cache_data__T_177_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_178_en & cache_data__T_178_mask) begin
      cache_data[cache_data__T_178_addr] <= cache_data__T_178_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_179_en & cache_data__T_179_mask) begin
      cache_data[cache_data__T_179_addr] <= cache_data__T_179_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_180_en & cache_data__T_180_mask) begin
      cache_data[cache_data__T_180_addr] <= cache_data__T_180_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_181_en & cache_data__T_181_mask) begin
      cache_data[cache_data__T_181_addr] <= cache_data__T_181_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_182_en & cache_data__T_182_mask) begin
      cache_data[cache_data__T_182_addr] <= cache_data__T_182_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_183_en & cache_data__T_183_mask) begin
      cache_data[cache_data__T_183_addr] <= cache_data__T_183_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_184_en & cache_data__T_184_mask) begin
      cache_data[cache_data__T_184_addr] <= cache_data__T_184_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_185_en & cache_data__T_185_mask) begin
      cache_data[cache_data__T_185_addr] <= cache_data__T_185_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_186_en & cache_data__T_186_mask) begin
      cache_data[cache_data__T_186_addr] <= cache_data__T_186_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_187_en & cache_data__T_187_mask) begin
      cache_data[cache_data__T_187_addr] <= cache_data__T_187_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_188_en & cache_data__T_188_mask) begin
      cache_data[cache_data__T_188_addr] <= cache_data__T_188_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_189_en & cache_data__T_189_mask) begin
      cache_data[cache_data__T_189_addr] <= cache_data__T_189_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_190_en & cache_data__T_190_mask) begin
      cache_data[cache_data__T_190_addr] <= cache_data__T_190_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_191_en & cache_data__T_191_mask) begin
      cache_data[cache_data__T_191_addr] <= cache_data__T_191_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_192_en & cache_data__T_192_mask) begin
      cache_data[cache_data__T_192_addr] <= cache_data__T_192_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_193_en & cache_data__T_193_mask) begin
      cache_data[cache_data__T_193_addr] <= cache_data__T_193_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_194_en & cache_data__T_194_mask) begin
      cache_data[cache_data__T_194_addr] <= cache_data__T_194_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_195_en & cache_data__T_195_mask) begin
      cache_data[cache_data__T_195_addr] <= cache_data__T_195_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_196_en & cache_data__T_196_mask) begin
      cache_data[cache_data__T_196_addr] <= cache_data__T_196_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_197_en & cache_data__T_197_mask) begin
      cache_data[cache_data__T_197_addr] <= cache_data__T_197_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_198_en & cache_data__T_198_mask) begin
      cache_data[cache_data__T_198_addr] <= cache_data__T_198_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_199_en & cache_data__T_199_mask) begin
      cache_data[cache_data__T_199_addr] <= cache_data__T_199_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_200_en & cache_data__T_200_mask) begin
      cache_data[cache_data__T_200_addr] <= cache_data__T_200_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_201_en & cache_data__T_201_mask) begin
      cache_data[cache_data__T_201_addr] <= cache_data__T_201_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_202_en & cache_data__T_202_mask) begin
      cache_data[cache_data__T_202_addr] <= cache_data__T_202_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_203_en & cache_data__T_203_mask) begin
      cache_data[cache_data__T_203_addr] <= cache_data__T_203_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_204_en & cache_data__T_204_mask) begin
      cache_data[cache_data__T_204_addr] <= cache_data__T_204_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_205_en & cache_data__T_205_mask) begin
      cache_data[cache_data__T_205_addr] <= cache_data__T_205_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_206_en & cache_data__T_206_mask) begin
      cache_data[cache_data__T_206_addr] <= cache_data__T_206_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_207_en & cache_data__T_207_mask) begin
      cache_data[cache_data__T_207_addr] <= cache_data__T_207_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_208_en & cache_data__T_208_mask) begin
      cache_data[cache_data__T_208_addr] <= cache_data__T_208_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_209_en & cache_data__T_209_mask) begin
      cache_data[cache_data__T_209_addr] <= cache_data__T_209_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_210_en & cache_data__T_210_mask) begin
      cache_data[cache_data__T_210_addr] <= cache_data__T_210_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_211_en & cache_data__T_211_mask) begin
      cache_data[cache_data__T_211_addr] <= cache_data__T_211_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_212_en & cache_data__T_212_mask) begin
      cache_data[cache_data__T_212_addr] <= cache_data__T_212_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_213_en & cache_data__T_213_mask) begin
      cache_data[cache_data__T_213_addr] <= cache_data__T_213_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_214_en & cache_data__T_214_mask) begin
      cache_data[cache_data__T_214_addr] <= cache_data__T_214_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_215_en & cache_data__T_215_mask) begin
      cache_data[cache_data__T_215_addr] <= cache_data__T_215_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_216_en & cache_data__T_216_mask) begin
      cache_data[cache_data__T_216_addr] <= cache_data__T_216_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_217_en & cache_data__T_217_mask) begin
      cache_data[cache_data__T_217_addr] <= cache_data__T_217_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_218_en & cache_data__T_218_mask) begin
      cache_data[cache_data__T_218_addr] <= cache_data__T_218_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_219_en & cache_data__T_219_mask) begin
      cache_data[cache_data__T_219_addr] <= cache_data__T_219_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_220_en & cache_data__T_220_mask) begin
      cache_data[cache_data__T_220_addr] <= cache_data__T_220_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_221_en & cache_data__T_221_mask) begin
      cache_data[cache_data__T_221_addr] <= cache_data__T_221_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_222_en & cache_data__T_222_mask) begin
      cache_data[cache_data__T_222_addr] <= cache_data__T_222_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_223_en & cache_data__T_223_mask) begin
      cache_data[cache_data__T_223_addr] <= cache_data__T_223_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_224_en & cache_data__T_224_mask) begin
      cache_data[cache_data__T_224_addr] <= cache_data__T_224_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_225_en & cache_data__T_225_mask) begin
      cache_data[cache_data__T_225_addr] <= cache_data__T_225_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_226_en & cache_data__T_226_mask) begin
      cache_data[cache_data__T_226_addr] <= cache_data__T_226_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_227_en & cache_data__T_227_mask) begin
      cache_data[cache_data__T_227_addr] <= cache_data__T_227_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_228_en & cache_data__T_228_mask) begin
      cache_data[cache_data__T_228_addr] <= cache_data__T_228_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_229_en & cache_data__T_229_mask) begin
      cache_data[cache_data__T_229_addr] <= cache_data__T_229_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_230_en & cache_data__T_230_mask) begin
      cache_data[cache_data__T_230_addr] <= cache_data__T_230_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_231_en & cache_data__T_231_mask) begin
      cache_data[cache_data__T_231_addr] <= cache_data__T_231_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_232_en & cache_data__T_232_mask) begin
      cache_data[cache_data__T_232_addr] <= cache_data__T_232_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_233_en & cache_data__T_233_mask) begin
      cache_data[cache_data__T_233_addr] <= cache_data__T_233_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_234_en & cache_data__T_234_mask) begin
      cache_data[cache_data__T_234_addr] <= cache_data__T_234_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_235_en & cache_data__T_235_mask) begin
      cache_data[cache_data__T_235_addr] <= cache_data__T_235_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_236_en & cache_data__T_236_mask) begin
      cache_data[cache_data__T_236_addr] <= cache_data__T_236_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_237_en & cache_data__T_237_mask) begin
      cache_data[cache_data__T_237_addr] <= cache_data__T_237_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_238_en & cache_data__T_238_mask) begin
      cache_data[cache_data__T_238_addr] <= cache_data__T_238_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_239_en & cache_data__T_239_mask) begin
      cache_data[cache_data__T_239_addr] <= cache_data__T_239_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_240_en & cache_data__T_240_mask) begin
      cache_data[cache_data__T_240_addr] <= cache_data__T_240_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_241_en & cache_data__T_241_mask) begin
      cache_data[cache_data__T_241_addr] <= cache_data__T_241_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_242_en & cache_data__T_242_mask) begin
      cache_data[cache_data__T_242_addr] <= cache_data__T_242_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_243_en & cache_data__T_243_mask) begin
      cache_data[cache_data__T_243_addr] <= cache_data__T_243_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_244_en & cache_data__T_244_mask) begin
      cache_data[cache_data__T_244_addr] <= cache_data__T_244_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_245_en & cache_data__T_245_mask) begin
      cache_data[cache_data__T_245_addr] <= cache_data__T_245_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_246_en & cache_data__T_246_mask) begin
      cache_data[cache_data__T_246_addr] <= cache_data__T_246_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_247_en & cache_data__T_247_mask) begin
      cache_data[cache_data__T_247_addr] <= cache_data__T_247_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_248_en & cache_data__T_248_mask) begin
      cache_data[cache_data__T_248_addr] <= cache_data__T_248_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_249_en & cache_data__T_249_mask) begin
      cache_data[cache_data__T_249_addr] <= cache_data__T_249_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_250_en & cache_data__T_250_mask) begin
      cache_data[cache_data__T_250_addr] <= cache_data__T_250_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_251_en & cache_data__T_251_mask) begin
      cache_data[cache_data__T_251_addr] <= cache_data__T_251_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_252_en & cache_data__T_252_mask) begin
      cache_data[cache_data__T_252_addr] <= cache_data__T_252_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_253_en & cache_data__T_253_mask) begin
      cache_data[cache_data__T_253_addr] <= cache_data__T_253_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_254_en & cache_data__T_254_mask) begin
      cache_data[cache_data__T_254_addr] <= cache_data__T_254_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_255_en & cache_data__T_255_mask) begin
      cache_data[cache_data__T_255_addr] <= cache_data__T_255_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_256_en & cache_data__T_256_mask) begin
      cache_data[cache_data__T_256_addr] <= cache_data__T_256_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_257_en & cache_data__T_257_mask) begin
      cache_data[cache_data__T_257_addr] <= cache_data__T_257_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_258_en & cache_data__T_258_mask) begin
      cache_data[cache_data__T_258_addr] <= cache_data__T_258_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_259_en & cache_data__T_259_mask) begin
      cache_data[cache_data__T_259_addr] <= cache_data__T_259_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_260_en & cache_data__T_260_mask) begin
      cache_data[cache_data__T_260_addr] <= cache_data__T_260_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_261_en & cache_data__T_261_mask) begin
      cache_data[cache_data__T_261_addr] <= cache_data__T_261_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_262_en & cache_data__T_262_mask) begin
      cache_data[cache_data__T_262_addr] <= cache_data__T_262_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_263_en & cache_data__T_263_mask) begin
      cache_data[cache_data__T_263_addr] <= cache_data__T_263_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_264_en & cache_data__T_264_mask) begin
      cache_data[cache_data__T_264_addr] <= cache_data__T_264_data; // @[icache.scala 91:18]
    end
    if(cache_data__T_265_en & cache_data__T_265_mask) begin
      cache_data[cache_data__T_265_addr] <= cache_data__T_265_data; // @[icache.scala 91:18]
    end
    if(cache_data_s1_entry_w_en & cache_data_s1_entry_w_mask) begin
      cache_data[cache_data_s1_entry_w_addr] <= cache_data_s1_entry_w_data; // @[icache.scala 91:18]
    end
    if (reset) begin
      s0_valid <= 1'h0;
    end else if (_T_273) begin
      s0_valid <= 1'h0;
    end else begin
      s0_valid <= _GEN_274;
    end
    if (reset) begin
      s0_in_is_cached <= 1'h0;
    end else if (_T_266) begin
      s0_in_is_cached <= io_in_req_bits_is_cached;
    end
    if (reset) begin
      s0_in_addr <= 32'h0;
    end else if (_T_266) begin
      s0_in_addr <= io_in_req_bits_addr;
    end
    if (reset) begin
      s0_in_len <= 2'h0;
    end else if (_T_266) begin
      s0_in_len <= 2'h3;
    end
    if (reset) begin
      s0_in_strb <= 4'h0;
    end else if (_T_266) begin
      s0_in_strb <= 4'hf;
    end
    if (reset) begin
      s1_in_addr <= 32'h0;
    end else if (s0_out_fire) begin
      s1_in_addr <= s0_in_addr;
    end
    if (reset) begin
      s1_valid <= 1'h0;
    end else if (_T_299) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= _GEN_283;
    end
    if (reset) begin
      s1_in_is_cached <= 1'h0;
    end else if (s0_out_fire) begin
      s1_in_is_cached <= s0_in_is_cached;
    end
    if (reset) begin
      s1_in_len <= 2'h0;
    end else if (s0_out_fire) begin
      s1_in_len <= s0_in_len;
    end
    if (reset) begin
      s1_in_strb <= 4'h0;
    end else if (s0_out_fire) begin
      s1_in_strb <= s0_in_strb;
    end
    if (reset) begin
      s1_req <= 1'h0;
    end else if (_T_309) begin
      s1_req <= 1'h0;
    end else begin
      s1_req <= _GEN_285;
    end
    if (reset) begin
      s1_resp <= 1'h0;
    end else if (_T_311) begin
      s1_resp <= 1'h0;
    end else begin
      s1_resp <= _GEN_287;
    end
    if (reset) begin
      s1_ex_wait <= 1'h0;
    end else if (_T_311) begin
      s1_ex_wait <= 1'h0;
    end else if (s1_ex_wait_en) begin
      s1_ex_wait <= io_ex_flush;
    end
  end
endmodule
module Divider(
  input         clock,
  input         reset,
  input         io_data_dividend_tvalid,
  input         io_data_divisor_tvalid,
  output        io_data_dout_tvalid,
  input  [39:0] io_data_dividend_tdata,
  input  [39:0] io_data_divisor_tdata,
  output [79:0] io_data_dout_tdata
);
  wire [40:0] quotient = $signed(io_data_dividend_tdata) / $signed(io_data_divisor_tdata); // @[top.scala 61:39]
  wire [39:0] remainder = $signed(io_data_dividend_tdata) % $signed(io_data_divisor_tdata); // @[top.scala 62:40]
  wire  _T_2 = io_data_dividend_tvalid & io_data_divisor_tvalid; // @[top.scala 65:43]
  wire [80:0] _T_3 = {quotient,remainder}; // @[Cat.scala 29:58]
  reg  pipePipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [79:0] pipePipe_bits; // @[Reg.scala 15:16]
  reg [95:0] _RAND_1;
  wire [80:0] _GEN_0 = _T_2 ? _T_3 : {{1'd0}, pipePipe_bits}; // @[Reg.scala 16:19]
  reg  pipePipe_valid_1; // @[Valid.scala 117:22]
  reg [31:0] _RAND_2;
  reg [79:0] pipePipe_bits_1; // @[Reg.scala 15:16]
  reg [95:0] _RAND_3;
  reg  pipePipe_valid_2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_4;
  reg [79:0] pipePipe_bits_2; // @[Reg.scala 15:16]
  reg [95:0] _RAND_5;
  reg  pipePipe_valid_3; // @[Valid.scala 117:22]
  reg [31:0] _RAND_6;
  reg [79:0] pipePipe_bits_3; // @[Reg.scala 15:16]
  reg [95:0] _RAND_7;
  reg  pipePipe_valid_4; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [79:0] pipePipe_bits_4; // @[Reg.scala 15:16]
  reg [95:0] _RAND_9;
  reg  pipePipe_valid_5; // @[Valid.scala 117:22]
  reg [31:0] _RAND_10;
  reg [79:0] pipePipe_bits_5; // @[Reg.scala 15:16]
  reg [95:0] _RAND_11;
  reg  pipePipe_valid_6; // @[Valid.scala 117:22]
  reg [31:0] _RAND_12;
  reg [79:0] pipePipe_bits_6; // @[Reg.scala 15:16]
  reg [95:0] _RAND_13;
  reg  pipePipe_valid_7; // @[Valid.scala 117:22]
  reg [31:0] _RAND_14;
  reg [79:0] pipePipe_bits_7; // @[Reg.scala 15:16]
  reg [95:0] _RAND_15;
  reg  pipePipe_valid_8; // @[Valid.scala 117:22]
  reg [31:0] _RAND_16;
  reg [79:0] pipePipe_bits_8; // @[Reg.scala 15:16]
  reg [95:0] _RAND_17;
  reg  pipePipe_valid_9; // @[Valid.scala 117:22]
  reg [31:0] _RAND_18;
  reg [79:0] pipePipe_bits_9; // @[Reg.scala 15:16]
  reg [95:0] _RAND_19;
  reg  pipePipe_valid_10; // @[Valid.scala 117:22]
  reg [31:0] _RAND_20;
  reg [79:0] pipePipe_bits_10; // @[Reg.scala 15:16]
  reg [95:0] _RAND_21;
  reg  pipePipe_valid_11; // @[Valid.scala 117:22]
  reg [31:0] _RAND_22;
  reg [79:0] pipePipe_bits_11; // @[Reg.scala 15:16]
  reg [95:0] _RAND_23;
  reg  pipePipe_valid_12; // @[Valid.scala 117:22]
  reg [31:0] _RAND_24;
  reg [79:0] pipePipe_bits_12; // @[Reg.scala 15:16]
  reg [95:0] _RAND_25;
  reg  pipePipe_valid_13; // @[Valid.scala 117:22]
  reg [31:0] _RAND_26;
  reg [79:0] pipePipe_bits_13; // @[Reg.scala 15:16]
  reg [95:0] _RAND_27;
  reg  pipePipe_valid_14; // @[Valid.scala 117:22]
  reg [31:0] _RAND_28;
  reg [79:0] pipePipe_bits_14; // @[Reg.scala 15:16]
  reg [95:0] _RAND_29;
  reg  pipePipe_valid_15; // @[Valid.scala 117:22]
  reg [31:0] _RAND_30;
  reg [79:0] pipePipe_bits_15; // @[Reg.scala 15:16]
  reg [95:0] _RAND_31;
  reg  pipePipe_valid_16; // @[Valid.scala 117:22]
  reg [31:0] _RAND_32;
  reg [79:0] pipePipe_bits_16; // @[Reg.scala 15:16]
  reg [95:0] _RAND_33;
  reg  pipePipe_valid_17; // @[Valid.scala 117:22]
  reg [31:0] _RAND_34;
  reg [79:0] pipePipe_bits_17; // @[Reg.scala 15:16]
  reg [95:0] _RAND_35;
  reg  pipePipe_valid_18; // @[Valid.scala 117:22]
  reg [31:0] _RAND_36;
  reg [79:0] pipePipe_bits_18; // @[Reg.scala 15:16]
  reg [95:0] _RAND_37;
  reg  pipePipe_valid_19; // @[Valid.scala 117:22]
  reg [31:0] _RAND_38;
  reg [79:0] pipePipe_bits_19; // @[Reg.scala 15:16]
  reg [95:0] _RAND_39;
  reg  pipePipe_valid_20; // @[Valid.scala 117:22]
  reg [31:0] _RAND_40;
  reg [79:0] pipePipe_bits_20; // @[Reg.scala 15:16]
  reg [95:0] _RAND_41;
  reg  pipePipe_valid_21; // @[Valid.scala 117:22]
  reg [31:0] _RAND_42;
  reg [79:0] pipePipe_bits_21; // @[Reg.scala 15:16]
  reg [95:0] _RAND_43;
  reg  pipePipe_valid_22; // @[Valid.scala 117:22]
  reg [31:0] _RAND_44;
  reg [79:0] pipePipe_bits_22; // @[Reg.scala 15:16]
  reg [95:0] _RAND_45;
  reg  pipePipe_valid_23; // @[Valid.scala 117:22]
  reg [31:0] _RAND_46;
  reg [79:0] pipePipe_bits_23; // @[Reg.scala 15:16]
  reg [95:0] _RAND_47;
  reg  pipePipe_valid_24; // @[Valid.scala 117:22]
  reg [31:0] _RAND_48;
  reg [79:0] pipePipe_bits_24; // @[Reg.scala 15:16]
  reg [95:0] _RAND_49;
  reg  pipePipe_valid_25; // @[Valid.scala 117:22]
  reg [31:0] _RAND_50;
  reg [79:0] pipePipe_bits_25; // @[Reg.scala 15:16]
  reg [95:0] _RAND_51;
  reg  pipePipe_valid_26; // @[Valid.scala 117:22]
  reg [31:0] _RAND_52;
  reg [79:0] pipePipe_bits_26; // @[Reg.scala 15:16]
  reg [95:0] _RAND_53;
  reg  pipePipe_valid_27; // @[Valid.scala 117:22]
  reg [31:0] _RAND_54;
  reg [79:0] pipePipe_bits_27; // @[Reg.scala 15:16]
  reg [95:0] _RAND_55;
  reg  pipePipe_valid_28; // @[Valid.scala 117:22]
  reg [31:0] _RAND_56;
  reg [79:0] pipePipe_bits_28; // @[Reg.scala 15:16]
  reg [95:0] _RAND_57;
  reg  pipePipe_valid_29; // @[Valid.scala 117:22]
  reg [31:0] _RAND_58;
  reg [79:0] pipePipe_bits_29; // @[Reg.scala 15:16]
  reg [95:0] _RAND_59;
  reg  pipePipe_valid_30; // @[Valid.scala 117:22]
  reg [31:0] _RAND_60;
  reg [79:0] pipePipe_bits_30; // @[Reg.scala 15:16]
  reg [95:0] _RAND_61;
  reg  pipePipe_valid_31; // @[Valid.scala 117:22]
  reg [31:0] _RAND_62;
  reg [79:0] pipePipe_bits_31; // @[Reg.scala 15:16]
  reg [95:0] _RAND_63;
  reg  pipePipe_valid_32; // @[Valid.scala 117:22]
  reg [31:0] _RAND_64;
  reg [79:0] pipePipe_bits_32; // @[Reg.scala 15:16]
  reg [95:0] _RAND_65;
  reg  pipePipe_valid_33; // @[Valid.scala 117:22]
  reg [31:0] _RAND_66;
  reg [79:0] pipePipe_bits_33; // @[Reg.scala 15:16]
  reg [95:0] _RAND_67;
  reg  pipePipe_valid_34; // @[Valid.scala 117:22]
  reg [31:0] _RAND_68;
  reg [79:0] pipePipe_bits_34; // @[Reg.scala 15:16]
  reg [95:0] _RAND_69;
  reg  pipePipe_valid_35; // @[Valid.scala 117:22]
  reg [31:0] _RAND_70;
  reg [79:0] pipePipe_bits_35; // @[Reg.scala 15:16]
  reg [95:0] _RAND_71;
  reg  pipePipe_valid_36; // @[Valid.scala 117:22]
  reg [31:0] _RAND_72;
  reg [79:0] pipePipe_bits_36; // @[Reg.scala 15:16]
  reg [95:0] _RAND_73;
  reg  pipePipe_valid_37; // @[Valid.scala 117:22]
  reg [31:0] _RAND_74;
  reg [79:0] pipePipe_bits_37; // @[Reg.scala 15:16]
  reg [95:0] _RAND_75;
  reg  pipePipe_valid_38; // @[Valid.scala 117:22]
  reg [31:0] _RAND_76;
  reg [79:0] pipePipe_bits_38; // @[Reg.scala 15:16]
  reg [95:0] _RAND_77;
  reg  pipePipe_valid_39; // @[Valid.scala 117:22]
  reg [31:0] _RAND_78;
  reg [79:0] pipePipe_bits_39; // @[Reg.scala 15:16]
  reg [95:0] _RAND_79;
  reg  pipePipe_valid_40; // @[Valid.scala 117:22]
  reg [31:0] _RAND_80;
  reg [79:0] pipePipe_bits_40; // @[Reg.scala 15:16]
  reg [95:0] _RAND_81;
  reg  pipePipe_valid_41; // @[Valid.scala 117:22]
  reg [31:0] _RAND_82;
  reg [79:0] pipePipe_bits_41; // @[Reg.scala 15:16]
  reg [95:0] _RAND_83;
  reg  pipePipe_valid_42; // @[Valid.scala 117:22]
  reg [31:0] _RAND_84;
  reg [79:0] pipePipe_bits_42; // @[Reg.scala 15:16]
  reg [95:0] _RAND_85;
  reg  pipePipe_valid_43; // @[Valid.scala 117:22]
  reg [31:0] _RAND_86;
  reg [79:0] pipePipe_bits_43; // @[Reg.scala 15:16]
  reg [95:0] _RAND_87;
  reg  pipePipe_valid_44; // @[Valid.scala 117:22]
  reg [31:0] _RAND_88;
  reg [79:0] pipePipe_bits_44; // @[Reg.scala 15:16]
  reg [95:0] _RAND_89;
  assign io_data_dout_tvalid = pipePipe_valid_44; // @[top.scala 70:23]
  assign io_data_dout_tdata = pipePipe_bits_44; // @[top.scala 71:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pipePipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  pipePipe_bits = _RAND_1[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  pipePipe_valid_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  pipePipe_bits_1 = _RAND_3[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  pipePipe_valid_2 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  pipePipe_bits_2 = _RAND_5[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  pipePipe_valid_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  pipePipe_bits_3 = _RAND_7[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  pipePipe_valid_4 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {3{`RANDOM}};
  pipePipe_bits_4 = _RAND_9[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  pipePipe_valid_5 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {3{`RANDOM}};
  pipePipe_bits_5 = _RAND_11[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  pipePipe_valid_6 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {3{`RANDOM}};
  pipePipe_bits_6 = _RAND_13[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  pipePipe_valid_7 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {3{`RANDOM}};
  pipePipe_bits_7 = _RAND_15[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  pipePipe_valid_8 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {3{`RANDOM}};
  pipePipe_bits_8 = _RAND_17[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  pipePipe_valid_9 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {3{`RANDOM}};
  pipePipe_bits_9 = _RAND_19[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  pipePipe_valid_10 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {3{`RANDOM}};
  pipePipe_bits_10 = _RAND_21[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  pipePipe_valid_11 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {3{`RANDOM}};
  pipePipe_bits_11 = _RAND_23[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  pipePipe_valid_12 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {3{`RANDOM}};
  pipePipe_bits_12 = _RAND_25[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  pipePipe_valid_13 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {3{`RANDOM}};
  pipePipe_bits_13 = _RAND_27[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  pipePipe_valid_14 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {3{`RANDOM}};
  pipePipe_bits_14 = _RAND_29[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  pipePipe_valid_15 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {3{`RANDOM}};
  pipePipe_bits_15 = _RAND_31[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  pipePipe_valid_16 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {3{`RANDOM}};
  pipePipe_bits_16 = _RAND_33[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  pipePipe_valid_17 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {3{`RANDOM}};
  pipePipe_bits_17 = _RAND_35[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  pipePipe_valid_18 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {3{`RANDOM}};
  pipePipe_bits_18 = _RAND_37[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  pipePipe_valid_19 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {3{`RANDOM}};
  pipePipe_bits_19 = _RAND_39[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  pipePipe_valid_20 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {3{`RANDOM}};
  pipePipe_bits_20 = _RAND_41[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  pipePipe_valid_21 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {3{`RANDOM}};
  pipePipe_bits_21 = _RAND_43[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  pipePipe_valid_22 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {3{`RANDOM}};
  pipePipe_bits_22 = _RAND_45[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  pipePipe_valid_23 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {3{`RANDOM}};
  pipePipe_bits_23 = _RAND_47[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  pipePipe_valid_24 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {3{`RANDOM}};
  pipePipe_bits_24 = _RAND_49[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  pipePipe_valid_25 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {3{`RANDOM}};
  pipePipe_bits_25 = _RAND_51[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  pipePipe_valid_26 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {3{`RANDOM}};
  pipePipe_bits_26 = _RAND_53[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  pipePipe_valid_27 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {3{`RANDOM}};
  pipePipe_bits_27 = _RAND_55[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  pipePipe_valid_28 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {3{`RANDOM}};
  pipePipe_bits_28 = _RAND_57[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  pipePipe_valid_29 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {3{`RANDOM}};
  pipePipe_bits_29 = _RAND_59[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  pipePipe_valid_30 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {3{`RANDOM}};
  pipePipe_bits_30 = _RAND_61[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  pipePipe_valid_31 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {3{`RANDOM}};
  pipePipe_bits_31 = _RAND_63[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  pipePipe_valid_32 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {3{`RANDOM}};
  pipePipe_bits_32 = _RAND_65[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  pipePipe_valid_33 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {3{`RANDOM}};
  pipePipe_bits_33 = _RAND_67[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  pipePipe_valid_34 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {3{`RANDOM}};
  pipePipe_bits_34 = _RAND_69[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  pipePipe_valid_35 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {3{`RANDOM}};
  pipePipe_bits_35 = _RAND_71[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  pipePipe_valid_36 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {3{`RANDOM}};
  pipePipe_bits_36 = _RAND_73[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  pipePipe_valid_37 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {3{`RANDOM}};
  pipePipe_bits_37 = _RAND_75[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  pipePipe_valid_38 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {3{`RANDOM}};
  pipePipe_bits_38 = _RAND_77[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  pipePipe_valid_39 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {3{`RANDOM}};
  pipePipe_bits_39 = _RAND_79[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  pipePipe_valid_40 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {3{`RANDOM}};
  pipePipe_bits_40 = _RAND_81[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  pipePipe_valid_41 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {3{`RANDOM}};
  pipePipe_bits_41 = _RAND_83[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  pipePipe_valid_42 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {3{`RANDOM}};
  pipePipe_bits_42 = _RAND_85[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  pipePipe_valid_43 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {3{`RANDOM}};
  pipePipe_bits_43 = _RAND_87[79:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  pipePipe_valid_44 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {3{`RANDOM}};
  pipePipe_bits_44 = _RAND_89[79:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pipePipe_valid <= 1'h0;
    end else begin
      pipePipe_valid <= _T_2;
    end
    pipePipe_bits <= _GEN_0[79:0];
    if (reset) begin
      pipePipe_valid_1 <= 1'h0;
    end else begin
      pipePipe_valid_1 <= pipePipe_valid;
    end
    if (pipePipe_valid) begin
      pipePipe_bits_1 <= pipePipe_bits;
    end
    if (reset) begin
      pipePipe_valid_2 <= 1'h0;
    end else begin
      pipePipe_valid_2 <= pipePipe_valid_1;
    end
    if (pipePipe_valid_1) begin
      pipePipe_bits_2 <= pipePipe_bits_1;
    end
    if (reset) begin
      pipePipe_valid_3 <= 1'h0;
    end else begin
      pipePipe_valid_3 <= pipePipe_valid_2;
    end
    if (pipePipe_valid_2) begin
      pipePipe_bits_3 <= pipePipe_bits_2;
    end
    if (reset) begin
      pipePipe_valid_4 <= 1'h0;
    end else begin
      pipePipe_valid_4 <= pipePipe_valid_3;
    end
    if (pipePipe_valid_3) begin
      pipePipe_bits_4 <= pipePipe_bits_3;
    end
    if (reset) begin
      pipePipe_valid_5 <= 1'h0;
    end else begin
      pipePipe_valid_5 <= pipePipe_valid_4;
    end
    if (pipePipe_valid_4) begin
      pipePipe_bits_5 <= pipePipe_bits_4;
    end
    if (reset) begin
      pipePipe_valid_6 <= 1'h0;
    end else begin
      pipePipe_valid_6 <= pipePipe_valid_5;
    end
    if (pipePipe_valid_5) begin
      pipePipe_bits_6 <= pipePipe_bits_5;
    end
    if (reset) begin
      pipePipe_valid_7 <= 1'h0;
    end else begin
      pipePipe_valid_7 <= pipePipe_valid_6;
    end
    if (pipePipe_valid_6) begin
      pipePipe_bits_7 <= pipePipe_bits_6;
    end
    if (reset) begin
      pipePipe_valid_8 <= 1'h0;
    end else begin
      pipePipe_valid_8 <= pipePipe_valid_7;
    end
    if (pipePipe_valid_7) begin
      pipePipe_bits_8 <= pipePipe_bits_7;
    end
    if (reset) begin
      pipePipe_valid_9 <= 1'h0;
    end else begin
      pipePipe_valid_9 <= pipePipe_valid_8;
    end
    if (pipePipe_valid_8) begin
      pipePipe_bits_9 <= pipePipe_bits_8;
    end
    if (reset) begin
      pipePipe_valid_10 <= 1'h0;
    end else begin
      pipePipe_valid_10 <= pipePipe_valid_9;
    end
    if (pipePipe_valid_9) begin
      pipePipe_bits_10 <= pipePipe_bits_9;
    end
    if (reset) begin
      pipePipe_valid_11 <= 1'h0;
    end else begin
      pipePipe_valid_11 <= pipePipe_valid_10;
    end
    if (pipePipe_valid_10) begin
      pipePipe_bits_11 <= pipePipe_bits_10;
    end
    if (reset) begin
      pipePipe_valid_12 <= 1'h0;
    end else begin
      pipePipe_valid_12 <= pipePipe_valid_11;
    end
    if (pipePipe_valid_11) begin
      pipePipe_bits_12 <= pipePipe_bits_11;
    end
    if (reset) begin
      pipePipe_valid_13 <= 1'h0;
    end else begin
      pipePipe_valid_13 <= pipePipe_valid_12;
    end
    if (pipePipe_valid_12) begin
      pipePipe_bits_13 <= pipePipe_bits_12;
    end
    if (reset) begin
      pipePipe_valid_14 <= 1'h0;
    end else begin
      pipePipe_valid_14 <= pipePipe_valid_13;
    end
    if (pipePipe_valid_13) begin
      pipePipe_bits_14 <= pipePipe_bits_13;
    end
    if (reset) begin
      pipePipe_valid_15 <= 1'h0;
    end else begin
      pipePipe_valid_15 <= pipePipe_valid_14;
    end
    if (pipePipe_valid_14) begin
      pipePipe_bits_15 <= pipePipe_bits_14;
    end
    if (reset) begin
      pipePipe_valid_16 <= 1'h0;
    end else begin
      pipePipe_valid_16 <= pipePipe_valid_15;
    end
    if (pipePipe_valid_15) begin
      pipePipe_bits_16 <= pipePipe_bits_15;
    end
    if (reset) begin
      pipePipe_valid_17 <= 1'h0;
    end else begin
      pipePipe_valid_17 <= pipePipe_valid_16;
    end
    if (pipePipe_valid_16) begin
      pipePipe_bits_17 <= pipePipe_bits_16;
    end
    if (reset) begin
      pipePipe_valid_18 <= 1'h0;
    end else begin
      pipePipe_valid_18 <= pipePipe_valid_17;
    end
    if (pipePipe_valid_17) begin
      pipePipe_bits_18 <= pipePipe_bits_17;
    end
    if (reset) begin
      pipePipe_valid_19 <= 1'h0;
    end else begin
      pipePipe_valid_19 <= pipePipe_valid_18;
    end
    if (pipePipe_valid_18) begin
      pipePipe_bits_19 <= pipePipe_bits_18;
    end
    if (reset) begin
      pipePipe_valid_20 <= 1'h0;
    end else begin
      pipePipe_valid_20 <= pipePipe_valid_19;
    end
    if (pipePipe_valid_19) begin
      pipePipe_bits_20 <= pipePipe_bits_19;
    end
    if (reset) begin
      pipePipe_valid_21 <= 1'h0;
    end else begin
      pipePipe_valid_21 <= pipePipe_valid_20;
    end
    if (pipePipe_valid_20) begin
      pipePipe_bits_21 <= pipePipe_bits_20;
    end
    if (reset) begin
      pipePipe_valid_22 <= 1'h0;
    end else begin
      pipePipe_valid_22 <= pipePipe_valid_21;
    end
    if (pipePipe_valid_21) begin
      pipePipe_bits_22 <= pipePipe_bits_21;
    end
    if (reset) begin
      pipePipe_valid_23 <= 1'h0;
    end else begin
      pipePipe_valid_23 <= pipePipe_valid_22;
    end
    if (pipePipe_valid_22) begin
      pipePipe_bits_23 <= pipePipe_bits_22;
    end
    if (reset) begin
      pipePipe_valid_24 <= 1'h0;
    end else begin
      pipePipe_valid_24 <= pipePipe_valid_23;
    end
    if (pipePipe_valid_23) begin
      pipePipe_bits_24 <= pipePipe_bits_23;
    end
    if (reset) begin
      pipePipe_valid_25 <= 1'h0;
    end else begin
      pipePipe_valid_25 <= pipePipe_valid_24;
    end
    if (pipePipe_valid_24) begin
      pipePipe_bits_25 <= pipePipe_bits_24;
    end
    if (reset) begin
      pipePipe_valid_26 <= 1'h0;
    end else begin
      pipePipe_valid_26 <= pipePipe_valid_25;
    end
    if (pipePipe_valid_25) begin
      pipePipe_bits_26 <= pipePipe_bits_25;
    end
    if (reset) begin
      pipePipe_valid_27 <= 1'h0;
    end else begin
      pipePipe_valid_27 <= pipePipe_valid_26;
    end
    if (pipePipe_valid_26) begin
      pipePipe_bits_27 <= pipePipe_bits_26;
    end
    if (reset) begin
      pipePipe_valid_28 <= 1'h0;
    end else begin
      pipePipe_valid_28 <= pipePipe_valid_27;
    end
    if (pipePipe_valid_27) begin
      pipePipe_bits_28 <= pipePipe_bits_27;
    end
    if (reset) begin
      pipePipe_valid_29 <= 1'h0;
    end else begin
      pipePipe_valid_29 <= pipePipe_valid_28;
    end
    if (pipePipe_valid_28) begin
      pipePipe_bits_29 <= pipePipe_bits_28;
    end
    if (reset) begin
      pipePipe_valid_30 <= 1'h0;
    end else begin
      pipePipe_valid_30 <= pipePipe_valid_29;
    end
    if (pipePipe_valid_29) begin
      pipePipe_bits_30 <= pipePipe_bits_29;
    end
    if (reset) begin
      pipePipe_valid_31 <= 1'h0;
    end else begin
      pipePipe_valid_31 <= pipePipe_valid_30;
    end
    if (pipePipe_valid_30) begin
      pipePipe_bits_31 <= pipePipe_bits_30;
    end
    if (reset) begin
      pipePipe_valid_32 <= 1'h0;
    end else begin
      pipePipe_valid_32 <= pipePipe_valid_31;
    end
    if (pipePipe_valid_31) begin
      pipePipe_bits_32 <= pipePipe_bits_31;
    end
    if (reset) begin
      pipePipe_valid_33 <= 1'h0;
    end else begin
      pipePipe_valid_33 <= pipePipe_valid_32;
    end
    if (pipePipe_valid_32) begin
      pipePipe_bits_33 <= pipePipe_bits_32;
    end
    if (reset) begin
      pipePipe_valid_34 <= 1'h0;
    end else begin
      pipePipe_valid_34 <= pipePipe_valid_33;
    end
    if (pipePipe_valid_33) begin
      pipePipe_bits_34 <= pipePipe_bits_33;
    end
    if (reset) begin
      pipePipe_valid_35 <= 1'h0;
    end else begin
      pipePipe_valid_35 <= pipePipe_valid_34;
    end
    if (pipePipe_valid_34) begin
      pipePipe_bits_35 <= pipePipe_bits_34;
    end
    if (reset) begin
      pipePipe_valid_36 <= 1'h0;
    end else begin
      pipePipe_valid_36 <= pipePipe_valid_35;
    end
    if (pipePipe_valid_35) begin
      pipePipe_bits_36 <= pipePipe_bits_35;
    end
    if (reset) begin
      pipePipe_valid_37 <= 1'h0;
    end else begin
      pipePipe_valid_37 <= pipePipe_valid_36;
    end
    if (pipePipe_valid_36) begin
      pipePipe_bits_37 <= pipePipe_bits_36;
    end
    if (reset) begin
      pipePipe_valid_38 <= 1'h0;
    end else begin
      pipePipe_valid_38 <= pipePipe_valid_37;
    end
    if (pipePipe_valid_37) begin
      pipePipe_bits_38 <= pipePipe_bits_37;
    end
    if (reset) begin
      pipePipe_valid_39 <= 1'h0;
    end else begin
      pipePipe_valid_39 <= pipePipe_valid_38;
    end
    if (pipePipe_valid_38) begin
      pipePipe_bits_39 <= pipePipe_bits_38;
    end
    if (reset) begin
      pipePipe_valid_40 <= 1'h0;
    end else begin
      pipePipe_valid_40 <= pipePipe_valid_39;
    end
    if (pipePipe_valid_39) begin
      pipePipe_bits_40 <= pipePipe_bits_39;
    end
    if (reset) begin
      pipePipe_valid_41 <= 1'h0;
    end else begin
      pipePipe_valid_41 <= pipePipe_valid_40;
    end
    if (pipePipe_valid_40) begin
      pipePipe_bits_41 <= pipePipe_bits_40;
    end
    if (reset) begin
      pipePipe_valid_42 <= 1'h0;
    end else begin
      pipePipe_valid_42 <= pipePipe_valid_41;
    end
    if (pipePipe_valid_41) begin
      pipePipe_bits_42 <= pipePipe_bits_41;
    end
    if (reset) begin
      pipePipe_valid_43 <= 1'h0;
    end else begin
      pipePipe_valid_43 <= pipePipe_valid_42;
    end
    if (pipePipe_valid_42) begin
      pipePipe_bits_43 <= pipePipe_bits_42;
    end
    if (reset) begin
      pipePipe_valid_44 <= 1'h0;
    end else begin
      pipePipe_valid_44 <= pipePipe_valid_43;
    end
    if (pipePipe_valid_43) begin
      pipePipe_bits_44 <= pipePipe_bits_43;
    end
  end
endmodule
module Multiplier(
  input         clock,
  input         reset,
  input  [32:0] io_data_a,
  input  [32:0] io_data_b,
  output [65:0] io_data_dout
);
  reg  pipePipe_valid; // @[Valid.scala 117:22]
  reg [31:0] _RAND_0;
  reg [65:0] pipePipe_bits; // @[Reg.scala 15:16]
  reg [95:0] _RAND_1;
  reg  pipePipe_valid_1; // @[Valid.scala 117:22]
  reg [31:0] _RAND_2;
  reg [65:0] pipePipe_bits_1; // @[Reg.scala 15:16]
  reg [95:0] _RAND_3;
  reg  pipePipe_valid_2; // @[Valid.scala 117:22]
  reg [31:0] _RAND_4;
  reg [65:0] pipePipe_bits_2; // @[Reg.scala 15:16]
  reg [95:0] _RAND_5;
  reg  pipePipe_valid_3; // @[Valid.scala 117:22]
  reg [31:0] _RAND_6;
  reg [65:0] pipePipe_bits_3; // @[Reg.scala 15:16]
  reg [95:0] _RAND_7;
  reg  pipePipe_valid_4; // @[Valid.scala 117:22]
  reg [31:0] _RAND_8;
  reg [65:0] pipePipe_bits_4; // @[Reg.scala 15:16]
  reg [95:0] _RAND_9;
  reg  pipePipe_valid_5; // @[Valid.scala 117:22]
  reg [31:0] _RAND_10;
  reg [65:0] pipePipe_bits_5; // @[Reg.scala 15:16]
  reg [95:0] _RAND_11;
  reg [65:0] pipePipe_bits_6; // @[Reg.scala 15:16]
  reg [95:0] _RAND_12;
  assign io_data_dout = pipePipe_bits_6; // @[top.scala 80:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pipePipe_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  pipePipe_bits = _RAND_1[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  pipePipe_valid_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {3{`RANDOM}};
  pipePipe_bits_1 = _RAND_3[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  pipePipe_valid_2 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {3{`RANDOM}};
  pipePipe_bits_2 = _RAND_5[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  pipePipe_valid_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {3{`RANDOM}};
  pipePipe_bits_3 = _RAND_7[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  pipePipe_valid_4 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {3{`RANDOM}};
  pipePipe_bits_4 = _RAND_9[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  pipePipe_valid_5 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {3{`RANDOM}};
  pipePipe_bits_5 = _RAND_11[65:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {3{`RANDOM}};
  pipePipe_bits_6 = _RAND_12[65:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pipePipe_valid <= 1'h0;
    end else begin
      pipePipe_valid <= 1'h1;
    end
    pipePipe_bits <= $signed(io_data_a) * $signed(io_data_b);
    if (reset) begin
      pipePipe_valid_1 <= 1'h0;
    end else begin
      pipePipe_valid_1 <= pipePipe_valid;
    end
    if (pipePipe_valid) begin
      pipePipe_bits_1 <= pipePipe_bits;
    end
    if (reset) begin
      pipePipe_valid_2 <= 1'h0;
    end else begin
      pipePipe_valid_2 <= pipePipe_valid_1;
    end
    if (pipePipe_valid_1) begin
      pipePipe_bits_2 <= pipePipe_bits_1;
    end
    if (reset) begin
      pipePipe_valid_3 <= 1'h0;
    end else begin
      pipePipe_valid_3 <= pipePipe_valid_2;
    end
    if (pipePipe_valid_2) begin
      pipePipe_bits_3 <= pipePipe_bits_2;
    end
    if (reset) begin
      pipePipe_valid_4 <= 1'h0;
    end else begin
      pipePipe_valid_4 <= pipePipe_valid_3;
    end
    if (pipePipe_valid_3) begin
      pipePipe_bits_4 <= pipePipe_bits_3;
    end
    if (reset) begin
      pipePipe_valid_5 <= 1'h0;
    end else begin
      pipePipe_valid_5 <= pipePipe_valid_4;
    end
    if (pipePipe_valid_4) begin
      pipePipe_bits_5 <= pipePipe_bits_4;
    end
    if (pipePipe_valid_5) begin
      pipePipe_bits_6 <= pipePipe_bits_5;
    end
  end
endmodule
module verilator_top(
  input         clock,
  input         reset,
  output        io_commit_valid,
  output [31:0] io_commit_pc,
  output [31:0] io_commit_instr,
  output        io_commit_ip7,
  output [31:0] io_commit_gpr_0,
  output [31:0] io_commit_gpr_1,
  output [31:0] io_commit_gpr_2,
  output [31:0] io_commit_gpr_3,
  output [31:0] io_commit_gpr_4,
  output [31:0] io_commit_gpr_5,
  output [31:0] io_commit_gpr_6,
  output [31:0] io_commit_gpr_7,
  output [31:0] io_commit_gpr_8,
  output [31:0] io_commit_gpr_9,
  output [31:0] io_commit_gpr_10,
  output [31:0] io_commit_gpr_11,
  output [31:0] io_commit_gpr_12,
  output [31:0] io_commit_gpr_13,
  output [31:0] io_commit_gpr_14,
  output [31:0] io_commit_gpr_15,
  output [31:0] io_commit_gpr_16,
  output [31:0] io_commit_gpr_17,
  output [31:0] io_commit_gpr_18,
  output [31:0] io_commit_gpr_19,
  output [31:0] io_commit_gpr_20,
  output [31:0] io_commit_gpr_21,
  output [31:0] io_commit_gpr_22,
  output [31:0] io_commit_gpr_23,
  output [31:0] io_commit_gpr_24,
  output [31:0] io_commit_gpr_25,
  output [31:0] io_commit_gpr_26,
  output [31:0] io_commit_gpr_27,
  output [31:0] io_commit_gpr_28,
  output [31:0] io_commit_gpr_29,
  output [31:0] io_commit_gpr_30,
  output [31:0] io_commit_gpr_31,
  output [4:0]  io_commit_rd_idx,
  output [31:0] io_commit_wdata,
  output        io_commit_wen,
  input         io_can_log_now
);
  wire  core_clock; // @[top.scala 89:20]
  wire  core_reset; // @[top.scala 89:20]
  wire  core_io_imem_req_ready; // @[top.scala 89:20]
  wire  core_io_imem_req_valid; // @[top.scala 89:20]
  wire  core_io_imem_req_bits_is_cached; // @[top.scala 89:20]
  wire [31:0] core_io_imem_req_bits_addr; // @[top.scala 89:20]
  wire  core_io_imem_resp_ready; // @[top.scala 89:20]
  wire  core_io_imem_resp_valid; // @[top.scala 89:20]
  wire [31:0] core_io_imem_resp_bits_data; // @[top.scala 89:20]
  wire  core_io_dmem_req_ready; // @[top.scala 89:20]
  wire  core_io_dmem_req_valid; // @[top.scala 89:20]
  wire  core_io_dmem_req_bits_is_cached; // @[top.scala 89:20]
  wire [31:0] core_io_dmem_req_bits_addr; // @[top.scala 89:20]
  wire [1:0] core_io_dmem_req_bits_len; // @[top.scala 89:20]
  wire [3:0] core_io_dmem_req_bits_strb; // @[top.scala 89:20]
  wire [31:0] core_io_dmem_req_bits_data; // @[top.scala 89:20]
  wire  core_io_dmem_req_bits_func; // @[top.scala 89:20]
  wire  core_io_dmem_resp_valid; // @[top.scala 89:20]
  wire [31:0] core_io_dmem_resp_bits_data; // @[top.scala 89:20]
  wire  core_io_icache_control_valid; // @[top.scala 89:20]
  wire [2:0] core_io_icache_control_bits_op; // @[top.scala 89:20]
  wire [31:0] core_io_icache_control_bits_addr; // @[top.scala 89:20]
  wire  core_io_commit_valid; // @[top.scala 89:20]
  wire [31:0] core_io_commit_pc; // @[top.scala 89:20]
  wire [31:0] core_io_commit_instr; // @[top.scala 89:20]
  wire  core_io_commit_ip7; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_0; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_1; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_2; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_3; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_4; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_5; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_6; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_7; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_8; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_9; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_10; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_11; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_12; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_13; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_14; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_15; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_16; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_17; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_18; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_19; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_20; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_21; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_22; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_23; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_24; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_25; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_26; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_27; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_28; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_29; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_30; // @[top.scala 89:20]
  wire [31:0] core_io_commit_gpr_31; // @[top.scala 89:20]
  wire [4:0] core_io_commit_rd_idx; // @[top.scala 89:20]
  wire [31:0] core_io_commit_wdata; // @[top.scala 89:20]
  wire  core_io_commit_wen; // @[top.scala 89:20]
  wire  core_io_br_flush; // @[top.scala 89:20]
  wire  core_io_ex_flush; // @[top.scala 89:20]
  wire [32:0] core_io_multiplier_data_a; // @[top.scala 89:20]
  wire [32:0] core_io_multiplier_data_b; // @[top.scala 89:20]
  wire [65:0] core_io_multiplier_data_dout; // @[top.scala 89:20]
  wire  core_io_divider_data_dividend_tvalid; // @[top.scala 89:20]
  wire  core_io_divider_data_divisor_tvalid; // @[top.scala 89:20]
  wire  core_io_divider_data_dout_tvalid; // @[top.scala 89:20]
  wire [39:0] core_io_divider_data_dividend_tdata; // @[top.scala 89:20]
  wire [39:0] core_io_divider_data_divisor_tdata; // @[top.scala 89:20]
  wire [79:0] core_io_divider_data_dout_tdata; // @[top.scala 89:20]
  wire  dev_clock; // @[top.scala 90:19]
  wire  dev_reset; // @[top.scala 90:19]
  wire  dev_in_req_ready; // @[top.scala 90:19]
  wire  dev_in_req_valid; // @[top.scala 90:19]
  wire  dev_in_req_bits_is_cached; // @[top.scala 90:19]
  wire [31:0] dev_in_req_bits_addr; // @[top.scala 90:19]
  wire [1:0] dev_in_req_bits_len; // @[top.scala 90:19]
  wire [3:0] dev_in_req_bits_strb; // @[top.scala 90:19]
  wire [31:0] dev_in_req_bits_data; // @[top.scala 90:19]
  wire  dev_in_req_bits_func; // @[top.scala 90:19]
  wire  dev_in_resp_ready; // @[top.scala 90:19]
  wire  dev_in_resp_valid; // @[top.scala 90:19]
  wire [31:0] dev_in_resp_bits_data; // @[top.scala 90:19]
  wire  crossbar_clock; // @[top.scala 91:24]
  wire  crossbar_reset; // @[top.scala 91:24]
  wire  crossbar_io_in_0_req_ready; // @[top.scala 91:24]
  wire  crossbar_io_in_0_req_valid; // @[top.scala 91:24]
  wire  crossbar_io_in_0_req_bits_is_cached; // @[top.scala 91:24]
  wire [31:0] crossbar_io_in_0_req_bits_addr; // @[top.scala 91:24]
  wire [1:0] crossbar_io_in_0_req_bits_len; // @[top.scala 91:24]
  wire [3:0] crossbar_io_in_0_req_bits_strb; // @[top.scala 91:24]
  wire  crossbar_io_in_0_resp_valid; // @[top.scala 91:24]
  wire [31:0] crossbar_io_in_0_resp_bits_data; // @[top.scala 91:24]
  wire  crossbar_io_in_1_req_ready; // @[top.scala 91:24]
  wire  crossbar_io_in_1_req_valid; // @[top.scala 91:24]
  wire  crossbar_io_in_1_req_bits_is_cached; // @[top.scala 91:24]
  wire [31:0] crossbar_io_in_1_req_bits_addr; // @[top.scala 91:24]
  wire [1:0] crossbar_io_in_1_req_bits_len; // @[top.scala 91:24]
  wire [3:0] crossbar_io_in_1_req_bits_strb; // @[top.scala 91:24]
  wire [31:0] crossbar_io_in_1_req_bits_data; // @[top.scala 91:24]
  wire  crossbar_io_in_1_req_bits_func; // @[top.scala 91:24]
  wire  crossbar_io_in_1_resp_valid; // @[top.scala 91:24]
  wire [31:0] crossbar_io_in_1_resp_bits_data; // @[top.scala 91:24]
  wire  crossbar_io_out_req_ready; // @[top.scala 91:24]
  wire  crossbar_io_out_req_valid; // @[top.scala 91:24]
  wire  crossbar_io_out_req_bits_is_cached; // @[top.scala 91:24]
  wire [31:0] crossbar_io_out_req_bits_addr; // @[top.scala 91:24]
  wire [1:0] crossbar_io_out_req_bits_len; // @[top.scala 91:24]
  wire [3:0] crossbar_io_out_req_bits_strb; // @[top.scala 91:24]
  wire [31:0] crossbar_io_out_req_bits_data; // @[top.scala 91:24]
  wire  crossbar_io_out_req_bits_func; // @[top.scala 91:24]
  wire  crossbar_io_out_resp_ready; // @[top.scala 91:24]
  wire  crossbar_io_out_resp_valid; // @[top.scala 91:24]
  wire [31:0] crossbar_io_out_resp_bits_data; // @[top.scala 91:24]
  wire  icache_clock; // @[top.scala 92:22]
  wire  icache_reset; // @[top.scala 92:22]
  wire  icache_io_in_req_ready; // @[top.scala 92:22]
  wire  icache_io_in_req_valid; // @[top.scala 92:22]
  wire  icache_io_in_req_bits_is_cached; // @[top.scala 92:22]
  wire [31:0] icache_io_in_req_bits_addr; // @[top.scala 92:22]
  wire  icache_io_in_resp_ready; // @[top.scala 92:22]
  wire  icache_io_in_resp_valid; // @[top.scala 92:22]
  wire [31:0] icache_io_in_resp_bits_data; // @[top.scala 92:22]
  wire  icache_io_out_req_ready; // @[top.scala 92:22]
  wire  icache_io_out_req_valid; // @[top.scala 92:22]
  wire  icache_io_out_req_bits_is_cached; // @[top.scala 92:22]
  wire [31:0] icache_io_out_req_bits_addr; // @[top.scala 92:22]
  wire [1:0] icache_io_out_req_bits_len; // @[top.scala 92:22]
  wire [3:0] icache_io_out_req_bits_strb; // @[top.scala 92:22]
  wire  icache_io_out_resp_ready; // @[top.scala 92:22]
  wire  icache_io_out_resp_valid; // @[top.scala 92:22]
  wire [31:0] icache_io_out_resp_bits_data; // @[top.scala 92:22]
  wire  icache_io_br_flush; // @[top.scala 92:22]
  wire  icache_io_ex_flush; // @[top.scala 92:22]
  wire  icache_io_control_valid; // @[top.scala 92:22]
  wire [2:0] icache_io_control_bits_op; // @[top.scala 92:22]
  wire [31:0] icache_io_control_bits_addr; // @[top.scala 92:22]
  wire  divider_clock; // @[top.scala 93:23]
  wire  divider_reset; // @[top.scala 93:23]
  wire  divider_io_data_dividend_tvalid; // @[top.scala 93:23]
  wire  divider_io_data_divisor_tvalid; // @[top.scala 93:23]
  wire  divider_io_data_dout_tvalid; // @[top.scala 93:23]
  wire [39:0] divider_io_data_dividend_tdata; // @[top.scala 93:23]
  wire [39:0] divider_io_data_divisor_tdata; // @[top.scala 93:23]
  wire [79:0] divider_io_data_dout_tdata; // @[top.scala 93:23]
  wire  multiplier_clock; // @[top.scala 94:26]
  wire  multiplier_reset; // @[top.scala 94:26]
  wire [32:0] multiplier_io_data_a; // @[top.scala 94:26]
  wire [32:0] multiplier_io_data_b; // @[top.scala 94:26]
  wire [65:0] multiplier_io_data_dout; // @[top.scala 94:26]
  Core core ( // @[top.scala 89:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_ready(core_io_imem_req_ready),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_is_cached(core_io_imem_req_bits_is_cached),
    .io_imem_req_bits_addr(core_io_imem_req_bits_addr),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_is_cached(core_io_dmem_req_bits_is_cached),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_len(core_io_dmem_req_bits_len),
    .io_dmem_req_bits_strb(core_io_dmem_req_bits_strb),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_req_bits_func(core_io_dmem_req_bits_func),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_icache_control_valid(core_io_icache_control_valid),
    .io_icache_control_bits_op(core_io_icache_control_bits_op),
    .io_icache_control_bits_addr(core_io_icache_control_bits_addr),
    .io_commit_valid(core_io_commit_valid),
    .io_commit_pc(core_io_commit_pc),
    .io_commit_instr(core_io_commit_instr),
    .io_commit_ip7(core_io_commit_ip7),
    .io_commit_gpr_0(core_io_commit_gpr_0),
    .io_commit_gpr_1(core_io_commit_gpr_1),
    .io_commit_gpr_2(core_io_commit_gpr_2),
    .io_commit_gpr_3(core_io_commit_gpr_3),
    .io_commit_gpr_4(core_io_commit_gpr_4),
    .io_commit_gpr_5(core_io_commit_gpr_5),
    .io_commit_gpr_6(core_io_commit_gpr_6),
    .io_commit_gpr_7(core_io_commit_gpr_7),
    .io_commit_gpr_8(core_io_commit_gpr_8),
    .io_commit_gpr_9(core_io_commit_gpr_9),
    .io_commit_gpr_10(core_io_commit_gpr_10),
    .io_commit_gpr_11(core_io_commit_gpr_11),
    .io_commit_gpr_12(core_io_commit_gpr_12),
    .io_commit_gpr_13(core_io_commit_gpr_13),
    .io_commit_gpr_14(core_io_commit_gpr_14),
    .io_commit_gpr_15(core_io_commit_gpr_15),
    .io_commit_gpr_16(core_io_commit_gpr_16),
    .io_commit_gpr_17(core_io_commit_gpr_17),
    .io_commit_gpr_18(core_io_commit_gpr_18),
    .io_commit_gpr_19(core_io_commit_gpr_19),
    .io_commit_gpr_20(core_io_commit_gpr_20),
    .io_commit_gpr_21(core_io_commit_gpr_21),
    .io_commit_gpr_22(core_io_commit_gpr_22),
    .io_commit_gpr_23(core_io_commit_gpr_23),
    .io_commit_gpr_24(core_io_commit_gpr_24),
    .io_commit_gpr_25(core_io_commit_gpr_25),
    .io_commit_gpr_26(core_io_commit_gpr_26),
    .io_commit_gpr_27(core_io_commit_gpr_27),
    .io_commit_gpr_28(core_io_commit_gpr_28),
    .io_commit_gpr_29(core_io_commit_gpr_29),
    .io_commit_gpr_30(core_io_commit_gpr_30),
    .io_commit_gpr_31(core_io_commit_gpr_31),
    .io_commit_rd_idx(core_io_commit_rd_idx),
    .io_commit_wdata(core_io_commit_wdata),
    .io_commit_wen(core_io_commit_wen),
    .io_br_flush(core_io_br_flush),
    .io_ex_flush(core_io_ex_flush),
    .io_multiplier_data_a(core_io_multiplier_data_a),
    .io_multiplier_data_b(core_io_multiplier_data_b),
    .io_multiplier_data_dout(core_io_multiplier_data_dout),
    .io_divider_data_dividend_tvalid(core_io_divider_data_dividend_tvalid),
    .io_divider_data_divisor_tvalid(core_io_divider_data_divisor_tvalid),
    .io_divider_data_dout_tvalid(core_io_divider_data_dout_tvalid),
    .io_divider_data_dividend_tdata(core_io_divider_data_dividend_tdata),
    .io_divider_data_divisor_tdata(core_io_divider_data_divisor_tdata),
    .io_divider_data_dout_tdata(core_io_divider_data_dout_tdata)
  );
  SimDev dev ( // @[top.scala 90:19]
    .clock(dev_clock),
    .reset(dev_reset),
    .in_req_ready(dev_in_req_ready),
    .in_req_valid(dev_in_req_valid),
    .in_req_bits_is_cached(dev_in_req_bits_is_cached),
    .in_req_bits_addr(dev_in_req_bits_addr),
    .in_req_bits_len(dev_in_req_bits_len),
    .in_req_bits_strb(dev_in_req_bits_strb),
    .in_req_bits_data(dev_in_req_bits_data),
    .in_req_bits_func(dev_in_req_bits_func),
    .in_resp_ready(dev_in_resp_ready),
    .in_resp_valid(dev_in_resp_valid),
    .in_resp_bits_data(dev_in_resp_bits_data)
  );
  CrossbarNx1 crossbar ( // @[top.scala 91:24]
    .clock(crossbar_clock),
    .reset(crossbar_reset),
    .io_in_0_req_ready(crossbar_io_in_0_req_ready),
    .io_in_0_req_valid(crossbar_io_in_0_req_valid),
    .io_in_0_req_bits_is_cached(crossbar_io_in_0_req_bits_is_cached),
    .io_in_0_req_bits_addr(crossbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_len(crossbar_io_in_0_req_bits_len),
    .io_in_0_req_bits_strb(crossbar_io_in_0_req_bits_strb),
    .io_in_0_resp_valid(crossbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_data(crossbar_io_in_0_resp_bits_data),
    .io_in_1_req_ready(crossbar_io_in_1_req_ready),
    .io_in_1_req_valid(crossbar_io_in_1_req_valid),
    .io_in_1_req_bits_is_cached(crossbar_io_in_1_req_bits_is_cached),
    .io_in_1_req_bits_addr(crossbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_len(crossbar_io_in_1_req_bits_len),
    .io_in_1_req_bits_strb(crossbar_io_in_1_req_bits_strb),
    .io_in_1_req_bits_data(crossbar_io_in_1_req_bits_data),
    .io_in_1_req_bits_func(crossbar_io_in_1_req_bits_func),
    .io_in_1_resp_valid(crossbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_data(crossbar_io_in_1_resp_bits_data),
    .io_out_req_ready(crossbar_io_out_req_ready),
    .io_out_req_valid(crossbar_io_out_req_valid),
    .io_out_req_bits_is_cached(crossbar_io_out_req_bits_is_cached),
    .io_out_req_bits_addr(crossbar_io_out_req_bits_addr),
    .io_out_req_bits_len(crossbar_io_out_req_bits_len),
    .io_out_req_bits_strb(crossbar_io_out_req_bits_strb),
    .io_out_req_bits_data(crossbar_io_out_req_bits_data),
    .io_out_req_bits_func(crossbar_io_out_req_bits_func),
    .io_out_resp_ready(crossbar_io_out_resp_ready),
    .io_out_resp_valid(crossbar_io_out_resp_valid),
    .io_out_resp_bits_data(crossbar_io_out_resp_bits_data)
  );
  SimICache icache ( // @[top.scala 92:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_in_req_ready(icache_io_in_req_ready),
    .io_in_req_valid(icache_io_in_req_valid),
    .io_in_req_bits_is_cached(icache_io_in_req_bits_is_cached),
    .io_in_req_bits_addr(icache_io_in_req_bits_addr),
    .io_in_resp_ready(icache_io_in_resp_ready),
    .io_in_resp_valid(icache_io_in_resp_valid),
    .io_in_resp_bits_data(icache_io_in_resp_bits_data),
    .io_out_req_ready(icache_io_out_req_ready),
    .io_out_req_valid(icache_io_out_req_valid),
    .io_out_req_bits_is_cached(icache_io_out_req_bits_is_cached),
    .io_out_req_bits_addr(icache_io_out_req_bits_addr),
    .io_out_req_bits_len(icache_io_out_req_bits_len),
    .io_out_req_bits_strb(icache_io_out_req_bits_strb),
    .io_out_resp_ready(icache_io_out_resp_ready),
    .io_out_resp_valid(icache_io_out_resp_valid),
    .io_out_resp_bits_data(icache_io_out_resp_bits_data),
    .io_br_flush(icache_io_br_flush),
    .io_ex_flush(icache_io_ex_flush),
    .io_control_valid(icache_io_control_valid),
    .io_control_bits_op(icache_io_control_bits_op),
    .io_control_bits_addr(icache_io_control_bits_addr)
  );
  Divider divider ( // @[top.scala 93:23]
    .clock(divider_clock),
    .reset(divider_reset),
    .io_data_dividend_tvalid(divider_io_data_dividend_tvalid),
    .io_data_divisor_tvalid(divider_io_data_divisor_tvalid),
    .io_data_dout_tvalid(divider_io_data_dout_tvalid),
    .io_data_dividend_tdata(divider_io_data_dividend_tdata),
    .io_data_divisor_tdata(divider_io_data_divisor_tdata),
    .io_data_dout_tdata(divider_io_data_dout_tdata)
  );
  Multiplier multiplier ( // @[top.scala 94:26]
    .clock(multiplier_clock),
    .reset(multiplier_reset),
    .io_data_a(multiplier_io_data_a),
    .io_data_b(multiplier_io_data_b),
    .io_data_dout(multiplier_io_data_dout)
  );
  assign io_commit_valid = core_io_commit_valid; // @[top.scala 120:18]
  assign io_commit_pc = core_io_commit_pc; // @[top.scala 120:18]
  assign io_commit_instr = core_io_commit_instr; // @[top.scala 120:18]
  assign io_commit_ip7 = core_io_commit_ip7; // @[top.scala 120:18]
  assign io_commit_gpr_0 = core_io_commit_gpr_0; // @[top.scala 120:18]
  assign io_commit_gpr_1 = core_io_commit_gpr_1; // @[top.scala 120:18]
  assign io_commit_gpr_2 = core_io_commit_gpr_2; // @[top.scala 120:18]
  assign io_commit_gpr_3 = core_io_commit_gpr_3; // @[top.scala 120:18]
  assign io_commit_gpr_4 = core_io_commit_gpr_4; // @[top.scala 120:18]
  assign io_commit_gpr_5 = core_io_commit_gpr_5; // @[top.scala 120:18]
  assign io_commit_gpr_6 = core_io_commit_gpr_6; // @[top.scala 120:18]
  assign io_commit_gpr_7 = core_io_commit_gpr_7; // @[top.scala 120:18]
  assign io_commit_gpr_8 = core_io_commit_gpr_8; // @[top.scala 120:18]
  assign io_commit_gpr_9 = core_io_commit_gpr_9; // @[top.scala 120:18]
  assign io_commit_gpr_10 = core_io_commit_gpr_10; // @[top.scala 120:18]
  assign io_commit_gpr_11 = core_io_commit_gpr_11; // @[top.scala 120:18]
  assign io_commit_gpr_12 = core_io_commit_gpr_12; // @[top.scala 120:18]
  assign io_commit_gpr_13 = core_io_commit_gpr_13; // @[top.scala 120:18]
  assign io_commit_gpr_14 = core_io_commit_gpr_14; // @[top.scala 120:18]
  assign io_commit_gpr_15 = core_io_commit_gpr_15; // @[top.scala 120:18]
  assign io_commit_gpr_16 = core_io_commit_gpr_16; // @[top.scala 120:18]
  assign io_commit_gpr_17 = core_io_commit_gpr_17; // @[top.scala 120:18]
  assign io_commit_gpr_18 = core_io_commit_gpr_18; // @[top.scala 120:18]
  assign io_commit_gpr_19 = core_io_commit_gpr_19; // @[top.scala 120:18]
  assign io_commit_gpr_20 = core_io_commit_gpr_20; // @[top.scala 120:18]
  assign io_commit_gpr_21 = core_io_commit_gpr_21; // @[top.scala 120:18]
  assign io_commit_gpr_22 = core_io_commit_gpr_22; // @[top.scala 120:18]
  assign io_commit_gpr_23 = core_io_commit_gpr_23; // @[top.scala 120:18]
  assign io_commit_gpr_24 = core_io_commit_gpr_24; // @[top.scala 120:18]
  assign io_commit_gpr_25 = core_io_commit_gpr_25; // @[top.scala 120:18]
  assign io_commit_gpr_26 = core_io_commit_gpr_26; // @[top.scala 120:18]
  assign io_commit_gpr_27 = core_io_commit_gpr_27; // @[top.scala 120:18]
  assign io_commit_gpr_28 = core_io_commit_gpr_28; // @[top.scala 120:18]
  assign io_commit_gpr_29 = core_io_commit_gpr_29; // @[top.scala 120:18]
  assign io_commit_gpr_30 = core_io_commit_gpr_30; // @[top.scala 120:18]
  assign io_commit_gpr_31 = core_io_commit_gpr_31; // @[top.scala 120:18]
  assign io_commit_rd_idx = core_io_commit_rd_idx; // @[top.scala 120:18]
  assign io_commit_wdata = core_io_commit_wdata; // @[top.scala 120:18]
  assign io_commit_wen = core_io_commit_wen; // @[top.scala 120:18]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_imem_req_ready = icache_io_in_req_ready; // @[top.scala 111:16]
  assign core_io_imem_resp_valid = icache_io_in_resp_valid; // @[top.scala 111:16]
  assign core_io_imem_resp_bits_data = icache_io_in_resp_bits_data; // @[top.scala 111:16]
  assign core_io_dmem_req_ready = crossbar_io_in_1_req_ready; // @[top.scala 114:17]
  assign core_io_dmem_resp_valid = crossbar_io_in_1_resp_valid; // @[top.scala 114:17]
  assign core_io_dmem_resp_bits_data = crossbar_io_in_1_resp_bits_data; // @[top.scala 114:17]
  assign core_io_multiplier_data_dout = multiplier_io_data_dout; // @[top.scala 109:17]
  assign core_io_divider_data_dout_tvalid = divider_io_data_dout_tvalid; // @[top.scala 108:14]
  assign core_io_divider_data_dout_tdata = divider_io_data_dout_tdata; // @[top.scala 108:14]
  assign dev_clock = clock; // @[top.scala 102:16]
  assign dev_reset = reset; // @[top.scala 103:16]
  assign dev_in_req_valid = crossbar_io_out_req_valid; // @[top.scala 118:19]
  assign dev_in_req_bits_is_cached = crossbar_io_out_req_bits_is_cached; // @[top.scala 118:19]
  assign dev_in_req_bits_addr = crossbar_io_out_req_bits_addr; // @[top.scala 118:19]
  assign dev_in_req_bits_len = crossbar_io_out_req_bits_len; // @[top.scala 118:19]
  assign dev_in_req_bits_strb = crossbar_io_out_req_bits_strb; // @[top.scala 118:19]
  assign dev_in_req_bits_data = crossbar_io_out_req_bits_data; // @[top.scala 118:19]
  assign dev_in_req_bits_func = crossbar_io_out_req_bits_func; // @[top.scala 118:19]
  assign dev_in_resp_ready = crossbar_io_out_resp_ready; // @[top.scala 118:19]
  assign crossbar_clock = clock;
  assign crossbar_reset = reset;
  assign crossbar_io_in_0_req_valid = icache_io_out_req_valid; // @[top.scala 113:17]
  assign crossbar_io_in_0_req_bits_is_cached = icache_io_out_req_bits_is_cached; // @[top.scala 113:17]
  assign crossbar_io_in_0_req_bits_addr = icache_io_out_req_bits_addr; // @[top.scala 113:17]
  assign crossbar_io_in_0_req_bits_len = icache_io_out_req_bits_len; // @[top.scala 113:17]
  assign crossbar_io_in_0_req_bits_strb = icache_io_out_req_bits_strb; // @[top.scala 113:17]
  assign crossbar_io_in_1_req_valid = core_io_dmem_req_valid; // @[top.scala 114:17]
  assign crossbar_io_in_1_req_bits_is_cached = core_io_dmem_req_bits_is_cached; // @[top.scala 114:17]
  assign crossbar_io_in_1_req_bits_addr = core_io_dmem_req_bits_addr; // @[top.scala 114:17]
  assign crossbar_io_in_1_req_bits_len = core_io_dmem_req_bits_len; // @[top.scala 114:17]
  assign crossbar_io_in_1_req_bits_strb = core_io_dmem_req_bits_strb; // @[top.scala 114:17]
  assign crossbar_io_in_1_req_bits_data = core_io_dmem_req_bits_data; // @[top.scala 114:17]
  assign crossbar_io_in_1_req_bits_func = core_io_dmem_req_bits_func; // @[top.scala 114:17]
  assign crossbar_io_out_req_ready = dev_in_req_ready; // @[top.scala 118:19]
  assign crossbar_io_out_resp_valid = dev_in_resp_valid; // @[top.scala 118:19]
  assign crossbar_io_out_resp_bits_data = dev_in_resp_bits_data; // @[top.scala 118:19]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_in_req_valid = core_io_imem_req_valid; // @[top.scala 111:16]
  assign icache_io_in_req_bits_is_cached = core_io_imem_req_bits_is_cached; // @[top.scala 111:16]
  assign icache_io_in_req_bits_addr = core_io_imem_req_bits_addr; // @[top.scala 111:16]
  assign icache_io_in_resp_ready = core_io_imem_resp_ready; // @[top.scala 111:16]
  assign icache_io_out_req_ready = crossbar_io_in_0_req_ready; // @[top.scala 113:17]
  assign icache_io_out_resp_valid = crossbar_io_in_0_resp_valid; // @[top.scala 113:17]
  assign icache_io_out_resp_bits_data = crossbar_io_in_0_resp_bits_data; // @[top.scala 113:17]
  assign icache_io_br_flush = core_io_br_flush; // @[top.scala 105:22]
  assign icache_io_ex_flush = core_io_ex_flush; // @[top.scala 106:22]
  assign icache_io_control_valid = core_io_icache_control_valid; // @[top.scala 116:21]
  assign icache_io_control_bits_op = core_io_icache_control_bits_op; // @[top.scala 116:21]
  assign icache_io_control_bits_addr = core_io_icache_control_bits_addr; // @[top.scala 116:21]
  assign divider_clock = clock;
  assign divider_reset = reset;
  assign divider_io_data_dividend_tvalid = core_io_divider_data_dividend_tvalid; // @[top.scala 108:14]
  assign divider_io_data_divisor_tvalid = core_io_divider_data_divisor_tvalid; // @[top.scala 108:14]
  assign divider_io_data_dividend_tdata = core_io_divider_data_dividend_tdata; // @[top.scala 108:14]
  assign divider_io_data_divisor_tdata = core_io_divider_data_divisor_tdata; // @[top.scala 108:14]
  assign multiplier_clock = clock;
  assign multiplier_reset = reset;
  assign multiplier_io_data_a = core_io_multiplier_data_a; // @[top.scala 109:17]
  assign multiplier_io_data_b = core_io_multiplier_data_b; // @[top.scala 109:17]
endmodule
